/******************************************************************************
 ** Logisim goes FPGA automatic generated Verilog code                       **
 **                                                                          **
 ** Component : RAM_DATA_RAM                                                 **
 **                                                                          **
 ******************************************************************************/

`timescale 1ns/1ps
module RAM_DATA_RAM( 
//                     displaySel,
//                     display,
                     addr,
                     clk,
                     d,
                     we,
                     q);

   /***************************************************************************
    ** Here the inputs are defined                                           **
    ***************************************************************************/
//   input [31:0] displaySel;
   input[13:0]  addr;
   input  clk;
   input[31:0]  d;
   input  we;
   

   /***************************************************************************
    ** Here the outputs are defined                                          **
    ***************************************************************************/
   output[31:0] q;
//   output [31:0] display;

	reg [31:0] mem[8740:0];
	always @ (posedge clk) begin
		if (we)
			mem[addr] <= d;
	end
	assign q = mem[addr];
//	assign q = displaySel[0] ? mem[10] :
//	                 displaySel[1] ? mem[11] :
//	                 displaySel[2] ? mem[12] :
//	                 displaySel[3] ? mem[13] :
//	                 displaySel[4] ? mem[14] :
//	                 displaySel[5] ? mem[15] :
//	                 displaySel[6] ? mem[16] :
//	                 displaySel[7] ? mem[17] :
//	                 displaySel[8] ? mem[18] :
//	                 displaySel[9] ? mem[19] :
//	                 displaySel[10] ? mem[20] :
//	                 displaySel[11] ? mem[30] :
//	                 displaySel[12] ? mem[100] :
//	                 displaySel[13] ? mem[300] :
//	                 displaySel[14] ? mem[500] :
//	                 displaySel[15] ? mem[700] : mem[addr];
	
	initial
    begin
        mem[14'd0] <= 32'hbf21257c;
        mem[14'd1] <= 32'h3f00e791;
        mem[14'd2] <= 32'h3e5bbb99;
        mem[14'd3] <= 32'hbecd0bf1;
        mem[14'd4] <= 32'h3a9eaefc;
        mem[14'd5] <= 32'h3ff89dda;
        mem[14'd6] <= 32'hbe33a817;
        mem[14'd7] <= 32'h3f837ba5;
        mem[14'd8] <= 32'hbffe9a26;
        mem[14'd9] <= 32'hbec6438e;
        mem[14'd900] <= 32'h3bace7e6;
        mem[14'd901] <= 32'hbc8b493f;
        mem[14'd902] <= 32'hbc701d60;
        mem[14'd903] <= 32'hbc8781a4;
        mem[14'd904] <= 32'hbb83864a;
        mem[14'd905] <= 32'hbc438158;
        mem[14'd906] <= 32'h3b93eb1a;
        mem[14'd907] <= 32'h3bdef518;
        mem[14'd908] <= 32'h3b94dcb2;
        mem[14'd909] <= 32'h3c476633;
        mem[14'd910] <= 32'h3a5b9564;
        mem[14'd911] <= 32'hbc8234e6;
        mem[14'd912] <= 32'hbc0e2867;
        mem[14'd913] <= 32'hba9602f4;
        mem[14'd914] <= 32'hbc99bb02;
        mem[14'd915] <= 32'h3708d930;
        mem[14'd916] <= 32'h3bf2dbbb;
        mem[14'd917] <= 32'hbac9f4b7;
        mem[14'd918] <= 32'hbc72873b;
        mem[14'd919] <= 32'hbc2a4712;
        mem[14'd920] <= 32'h3c26c5b4;
        mem[14'd921] <= 32'hbc36b8d9;
        mem[14'd922] <= 32'h3cb3de6e;
        mem[14'd923] <= 32'hbc49839e;
        mem[14'd924] <= 32'h3c277dd4;
        mem[14'd925] <= 32'h38c120d1;
        mem[14'd926] <= 32'h3bb5d50f;
        mem[14'd927] <= 32'h3c8fe462;
        mem[14'd928] <= 32'hbc7d75e9;
        mem[14'd929] <= 32'h3bae5cf3;
        mem[14'd930] <= 32'hbb45333c;
        mem[14'd931] <= 32'h39c099f8;
        mem[14'd932] <= 32'hb9b81cd6;
        mem[14'd933] <= 32'h3b8da84a;
        mem[14'd934] <= 32'hbb7b848a;
        mem[14'd935] <= 32'hbc266cf1;
        mem[14'd936] <= 32'h3abeadef;
        mem[14'd937] <= 32'h3b47fab1;
        mem[14'd938] <= 32'h3c184a88;
        mem[14'd939] <= 32'h3c8855f2;
        mem[14'd940] <= 32'h3cbf4a68;
        mem[14'd941] <= 32'h3c5f9a2d;
        mem[14'd942] <= 32'hbb6c4db9;
        mem[14'd943] <= 32'hbbb8d535;
        mem[14'd944] <= 32'h3d0233eb;
        mem[14'd945] <= 32'h3c80fb80;
        mem[14'd946] <= 32'h3a434b70;
        mem[14'd947] <= 32'h3c87dbbe;
        mem[14'd948] <= 32'hbba5b80f;
        mem[14'd949] <= 32'h3c0f9821;
        mem[14'd950] <= 32'h3b9f2b08;
        mem[14'd951] <= 32'h3cb53231;
        mem[14'd952] <= 32'hbc09e18b;
        mem[14'd953] <= 32'h3acf131d;
        mem[14'd954] <= 32'h3b87d6b4;
        mem[14'd955] <= 32'h3b42d73c;
        mem[14'd956] <= 32'h3c5340c0;
        mem[14'd957] <= 32'h3b45184a;
        mem[14'd958] <= 32'hb9919274;
        mem[14'd959] <= 32'h3c1d8304;
        mem[14'd960] <= 32'hbb9aab33;
        mem[14'd961] <= 32'h3bd76a97;
        mem[14'd962] <= 32'hbba16b10;
        mem[14'd963] <= 32'hbc3771bf;
        mem[14'd964] <= 32'hbc09346f;
        mem[14'd965] <= 32'hbb4f7bb5;
        mem[14'd966] <= 32'hbc926435;
        mem[14'd967] <= 32'hbc889e4e;
        mem[14'd968] <= 32'hbcc924c2;
        mem[14'd969] <= 32'hbd051a4e;
        mem[14'd970] <= 32'hbda3e9e7;
        mem[14'd971] <= 32'hbdb126f4;
        mem[14'd972] <= 32'hbd722cf6;
        mem[14'd973] <= 32'hbcdb1d1e;
        mem[14'd974] <= 32'hbcc320b4;
        mem[14'd975] <= 32'hbc1b4ac7;
        mem[14'd976] <= 32'hbd044c9c;
        mem[14'd977] <= 32'hbb9dc383;
        mem[14'd978] <= 32'hbb2269e0;
        mem[14'd979] <= 32'hbc125a0c;
        mem[14'd980] <= 32'hbc734687;
        mem[14'd981] <= 32'h3ac895cc;
        mem[14'd982] <= 32'h3c5608fe;
        mem[14'd983] <= 32'hbbbf7694;
        mem[14'd984] <= 32'hbbfcbc62;
        mem[14'd985] <= 32'hbbee3e69;
        mem[14'd986] <= 32'hbca05300;
        mem[14'd987] <= 32'h3c988d86;
        mem[14'd988] <= 32'hbb012ff6;
        mem[14'd989] <= 32'hbcd56a53;
        mem[14'd990] <= 32'hbceb6f2f;
        mem[14'd991] <= 32'hbd3b91cf;
        mem[14'd992] <= 32'h3a978717;
        mem[14'd993] <= 32'hbd49f83f;
        mem[14'd994] <= 32'hbcf81b46;
        mem[14'd995] <= 32'hbbf01393;
        mem[14'd996] <= 32'hbd0771b1;
        mem[14'd997] <= 32'h3c3d786f;
        mem[14'd998] <= 32'h3cbae9b8;
        mem[14'd999] <= 32'hbcbab230;
        mem[14'd1000] <= 32'hbcc8b677;
        mem[14'd1001] <= 32'hbccf239a;
        mem[14'd1002] <= 32'hbe1225c5;
        mem[14'd1003] <= 32'hbe13a7b2;
        mem[14'd1004] <= 32'hbdf136b0;
        mem[14'd1005] <= 32'hbdcb472b;
        mem[14'd1006] <= 32'hbd86cdb4;
        mem[14'd1007] <= 32'hbc9fbf21;
        mem[14'd1008] <= 32'hbcdaedd5;
        mem[14'd1009] <= 32'h3bde4927;
        mem[14'd1010] <= 32'h3a2fe0a7;
        mem[14'd1011] <= 32'hbc0490e3;
        mem[14'd1012] <= 32'hbb463024;
        mem[14'd1013] <= 32'h3c692ef4;
        mem[14'd1014] <= 32'hbb84b610;
        mem[14'd1015] <= 32'hbbbb870d;
        mem[14'd1016] <= 32'hbbacf466;
        mem[14'd1017] <= 32'hbd0128d8;
        mem[14'd1018] <= 32'hbd47f7ee;
        mem[14'd1019] <= 32'hbcfc1dd6;
        mem[14'd1020] <= 32'h3c4fd765;
        mem[14'd1021] <= 32'h3d0d61db;
        mem[14'd1022] <= 32'h3b75d6ba;
        mem[14'd1023] <= 32'h3d3363c4;
        mem[14'd1024] <= 32'hbc311390;
        mem[14'd1025] <= 32'h3cfae724;
        mem[14'd1026] <= 32'hbcb199fe;
        mem[14'd1027] <= 32'h3d17fad7;
        mem[14'd1028] <= 32'hbc8c3b85;
        mem[14'd1029] <= 32'h3d5c5af4;
        mem[14'd1030] <= 32'hbd1b9e9a;
        mem[14'd1031] <= 32'hbdca7104;
        mem[14'd1032] <= 32'hbdbd4bd4;
        mem[14'd1033] <= 32'hbdbf32ff;
        mem[14'd1034] <= 32'hbdce5d1b;
        mem[14'd1035] <= 32'hbd6df165;
        mem[14'd1036] <= 32'hbd94b5ef;
        mem[14'd1037] <= 32'hbcabdf23;
        mem[14'd1038] <= 32'hb9b78231;
        mem[14'd1039] <= 32'h3b12431c;
        mem[14'd1040] <= 32'hbbbf0709;
        mem[14'd1041] <= 32'h3b1892b2;
        mem[14'd1042] <= 32'hbb3c1f64;
        mem[14'd1043] <= 32'h3bce1571;
        mem[14'd1044] <= 32'hbc8f3e96;
        mem[14'd1045] <= 32'hbd981c6a;
        mem[14'd1046] <= 32'hbd08a0ea;
        mem[14'd1047] <= 32'hbcc60966;
        mem[14'd1048] <= 32'hbb7bfd4b;
        mem[14'd1049] <= 32'h3c88b800;
        mem[14'd1050] <= 32'h3dd16dfc;
        mem[14'd1051] <= 32'h3d7d47f9;
        mem[14'd1052] <= 32'h3bb0b0ab;
        mem[14'd1053] <= 32'h3e2b7458;
        mem[14'd1054] <= 32'h3e5c8450;
        mem[14'd1055] <= 32'h3e2a774e;
        mem[14'd1056] <= 32'h3e188678;
        mem[14'd1057] <= 32'h3e731214;
        mem[14'd1058] <= 32'h3e5f8064;
        mem[14'd1059] <= 32'h3d863aba;
        mem[14'd1060] <= 32'hbccaec70;
        mem[14'd1061] <= 32'h3cc16e78;
        mem[14'd1062] <= 32'hbc674308;
        mem[14'd1063] <= 32'hbdf6f3d3;
        mem[14'd1064] <= 32'hbde8e089;
        mem[14'd1065] <= 32'hbd87a7cb;
        mem[14'd1066] <= 32'hbcb7210e;
        mem[14'd1067] <= 32'h3c0d0542;
        mem[14'd1068] <= 32'hbb6365c5;
        mem[14'd1069] <= 32'h3c62e1bd;
        mem[14'd1070] <= 32'hbb113753;
        mem[14'd1071] <= 32'hbbc75117;
        mem[14'd1072] <= 32'hbd1e62bd;
        mem[14'd1073] <= 32'hbd22ea00;
        mem[14'd1074] <= 32'hbcce2039;
        mem[14'd1075] <= 32'hbca7350f;
        mem[14'd1076] <= 32'hbd4144f8;
        mem[14'd1077] <= 32'hbdc60501;
        mem[14'd1078] <= 32'h3cf7e2dc;
        mem[14'd1079] <= 32'h3c2804ff;
        mem[14'd1080] <= 32'hbcd586a9;
        mem[14'd1081] <= 32'h3e273592;
        mem[14'd1082] <= 32'h3e1d2322;
        mem[14'd1083] <= 32'h3d418fc3;
        mem[14'd1084] <= 32'h3e07387f;
        mem[14'd1085] <= 32'h3e58c931;
        mem[14'd1086] <= 32'h3e814c41;
        mem[14'd1087] <= 32'h3e0ec8c8;
        mem[14'd1088] <= 32'h3da24cc4;
        mem[14'd1089] <= 32'h3e503ba8;
        mem[14'd1090] <= 32'h3e4b5014;
        mem[14'd1091] <= 32'hbcd788f7;
        mem[14'd1092] <= 32'hbe523fcd;
        mem[14'd1093] <= 32'hbe2dadba;
        mem[14'd1094] <= 32'hbd2dd304;
        mem[14'd1095] <= 32'hbc4aaad4;
        mem[14'd1096] <= 32'hbc4c163c;
        mem[14'd1097] <= 32'hbade937d;
        mem[14'd1098] <= 32'hbc21ef0a;
        mem[14'd1099] <= 32'hbbab16f8;
        mem[14'd1100] <= 32'hbd1e3ee7;
        mem[14'd1101] <= 32'hbd55ba04;
        mem[14'd1102] <= 32'hbcaa55cf;
        mem[14'd1103] <= 32'hbd495b6f;
        mem[14'd1104] <= 32'hbe0e833b;
        mem[14'd1105] <= 32'h3ba2931b;
        mem[14'd1106] <= 32'h3d6a10d4;
        mem[14'd1107] <= 32'h3d95a0ea;
        mem[14'd1108] <= 32'h3cbfdf76;
        mem[14'd1109] <= 32'h3df639a4;
        mem[14'd1110] <= 32'h3dc246ff;
        mem[14'd1111] <= 32'h3d88c765;
        mem[14'd1112] <= 32'h3db9c930;
        mem[14'd1113] <= 32'h3e82b736;
        mem[14'd1114] <= 32'h3e65a007;
        mem[14'd1115] <= 32'h3e246541;
        mem[14'd1116] <= 32'h3d4c0493;
        mem[14'd1117] <= 32'h3d88bebc;
        mem[14'd1118] <= 32'h3e0df3b2;
        mem[14'd1119] <= 32'h3e0e7c7e;
        mem[14'd1120] <= 32'hbdc1b72f;
        mem[14'd1121] <= 32'hbe408285;
        mem[14'd1122] <= 32'hbd8cdbef;
        mem[14'd1123] <= 32'hbb224b97;
        mem[14'd1124] <= 32'h3c069751;
        mem[14'd1125] <= 32'h3b602b93;
        mem[14'd1126] <= 32'h3bc9a86e;
        mem[14'd1127] <= 32'hbc5911d6;
        mem[14'd1128] <= 32'hbd828b94;
        mem[14'd1129] <= 32'hbd74647e;
        mem[14'd1130] <= 32'hbd7c4474;
        mem[14'd1131] <= 32'hbd918ec0;
        mem[14'd1132] <= 32'hbd72d020;
        mem[14'd1133] <= 32'h3d8e9cf6;
        mem[14'd1134] <= 32'h3d8d9b27;
        mem[14'd1135] <= 32'h3bfe894f;
        mem[14'd1136] <= 32'h3dbc2677;
        mem[14'd1137] <= 32'h3d26e5ba;
        mem[14'd1138] <= 32'h3e32fba2;
        mem[14'd1139] <= 32'h3e62e666;
        mem[14'd1140] <= 32'h3ec4fbc1;
        mem[14'd1141] <= 32'h3e9337dc;
        mem[14'd1142] <= 32'h3e592555;
        mem[14'd1143] <= 32'h3db7531d;
        mem[14'd1144] <= 32'h3d873383;
        mem[14'd1145] <= 32'h3d78728b;
        mem[14'd1146] <= 32'h3e413575;
        mem[14'd1147] <= 32'h3e98f7ab;
        mem[14'd1148] <= 32'h3d1c386e;
        mem[14'd1149] <= 32'hbe38dc2f;
        mem[14'd1150] <= 32'hbd5d023b;
        mem[14'd1151] <= 32'h3bec76cc;
        mem[14'd1152] <= 32'hbbd78046;
        mem[14'd1153] <= 32'h3acdfee4;
        mem[14'd1154] <= 32'hba90d73c;
        mem[14'd1155] <= 32'hbc9364fb;
        mem[14'd1156] <= 32'hbd656e24;
        mem[14'd1157] <= 32'hbd272dc4;
        mem[14'd1158] <= 32'hbd92535e;
        mem[14'd1159] <= 32'hbdb10c32;
        mem[14'd1160] <= 32'hbdc111f8;
        mem[14'd1161] <= 32'h3c89f916;
        mem[14'd1162] <= 32'h3da38797;
        mem[14'd1163] <= 32'hbce2c72e;
        mem[14'd1164] <= 32'h3d3e0343;
        mem[14'd1165] <= 32'h3e4622c5;
        mem[14'd1166] <= 32'h3d9c5e6d;
        mem[14'd1167] <= 32'hbc953f8d;
        mem[14'd1168] <= 32'h3e22b314;
        mem[14'd1169] <= 32'h3e8fc753;
        mem[14'd1170] <= 32'h3e8230b7;
        mem[14'd1171] <= 32'h3e6fe464;
        mem[14'd1172] <= 32'h3df6a08a;
        mem[14'd1173] <= 32'hbc87c99c;
        mem[14'd1174] <= 32'h3de9eeed;
        mem[14'd1175] <= 32'h3eb2a273;
        mem[14'd1176] <= 32'h3e0d1a96;
        mem[14'd1177] <= 32'hbe3bf841;
        mem[14'd1178] <= 32'hbd37e4e4;
        mem[14'd1179] <= 32'h3c8ea289;
        mem[14'd1180] <= 32'hbc2aaaa8;
        mem[14'd1181] <= 32'h3bfcb565;
        mem[14'd1182] <= 32'h3c0351b6;
        mem[14'd1183] <= 32'hbc52bc46;
        mem[14'd1184] <= 32'hbd618f41;
        mem[14'd1185] <= 32'hbd075e3d;
        mem[14'd1186] <= 32'hbd9b2dbf;
        mem[14'd1187] <= 32'hbd9cdf44;
        mem[14'd1188] <= 32'hbd036216;
        mem[14'd1189] <= 32'h3d3aedad;
        mem[14'd1190] <= 32'hbda985e4;
        mem[14'd1191] <= 32'h3cc3484d;
        mem[14'd1192] <= 32'h3cda6b58;
        mem[14'd1193] <= 32'h3da62b2d;
        mem[14'd1194] <= 32'h3acd882f;
        mem[14'd1195] <= 32'hbe0fd47d;
        mem[14'd1196] <= 32'hbccd8d3e;
        mem[14'd1197] <= 32'h3e75ae4b;
        mem[14'd1198] <= 32'h3e6f125b;
        mem[14'd1199] <= 32'h3dc22a0c;
        mem[14'd1200] <= 32'h3e0e8aa7;
        mem[14'd1201] <= 32'h3db8d0dc;
        mem[14'd1202] <= 32'h3e5f39d3;
        mem[14'd1203] <= 32'h3ebf0a53;
        mem[14'd1204] <= 32'h3e59b845;
        mem[14'd1205] <= 32'hbe235e9b;
        mem[14'd1206] <= 32'hbd823115;
        mem[14'd1207] <= 32'hbc33c741;
        mem[14'd1208] <= 32'h3bc0714a;
        mem[14'd1209] <= 32'hbb528221;
        mem[14'd1210] <= 32'h3be4d8bd;
        mem[14'd1211] <= 32'h3b064f23;
        mem[14'd1212] <= 32'hbdd23ba2;
        mem[14'd1213] <= 32'hbdd0950b;
        mem[14'd1214] <= 32'h3bb63df5;
        mem[14'd1215] <= 32'h3ce483ad;
        mem[14'd1216] <= 32'hbc1926f4;
        mem[14'd1217] <= 32'hbdc750df;
        mem[14'd1218] <= 32'hbd8c4a45;
        mem[14'd1219] <= 32'hbc236a0a;
        mem[14'd1220] <= 32'hbdc917a3;
        mem[14'd1221] <= 32'hbd80b4be;
        mem[14'd1222] <= 32'hbeac78f4;
        mem[14'd1223] <= 32'hbf0a663f;
        mem[14'd1224] <= 32'hbef3196f;
        mem[14'd1225] <= 32'hbd71e930;
        mem[14'd1226] <= 32'hbd1ff1bc;
        mem[14'd1227] <= 32'h3dabef12;
        mem[14'd1228] <= 32'h3e200256;
        mem[14'd1229] <= 32'h3e67edc9;
        mem[14'd1230] <= 32'h3e6b21f5;
        mem[14'd1231] <= 32'h3ea7955c;
        mem[14'd1232] <= 32'h3e85a2e7;
        mem[14'd1233] <= 32'hbdb85a0a;
        mem[14'd1234] <= 32'hbd2b38be;
        mem[14'd1235] <= 32'hbc39d6a6;
        mem[14'd1236] <= 32'h3bd9198a;
        mem[14'd1237] <= 32'hbc654cd9;
        mem[14'd1238] <= 32'hbbe3a912;
        mem[14'd1239] <= 32'hbcaf2a84;
        mem[14'd1240] <= 32'hbdc2e430;
        mem[14'd1241] <= 32'hbca7a4bb;
        mem[14'd1242] <= 32'h3e1057e8;
        mem[14'd1243] <= 32'h3d5f4a37;
        mem[14'd1244] <= 32'hbc6b1b3e;
        mem[14'd1245] <= 32'hbc86188b;
        mem[14'd1246] <= 32'h3ce30868;
        mem[14'd1247] <= 32'h3bfb8706;
        mem[14'd1248] <= 32'h3d9660d1;
        mem[14'd1249] <= 32'hbd92620f;
        mem[14'd1250] <= 32'hbeff21d1;
        mem[14'd1251] <= 32'hbf36a9b8;
        mem[14'd1252] <= 32'hbf16e19e;
        mem[14'd1253] <= 32'hbe2f9451;
        mem[14'd1254] <= 32'hbd1acd1e;
        mem[14'd1255] <= 32'h3d465d1e;
        mem[14'd1256] <= 32'h3d558672;
        mem[14'd1257] <= 32'h3e03c497;
        mem[14'd1258] <= 32'h3e9230c7;
        mem[14'd1259] <= 32'h3ec4c108;
        mem[14'd1260] <= 32'h3eb5eef5;
        mem[14'd1261] <= 32'hbbed91f3;
        mem[14'd1262] <= 32'hbcb1d260;
        mem[14'd1263] <= 32'h3bb7385b;
        mem[14'd1264] <= 32'hbc4ccb29;
        mem[14'd1265] <= 32'hbab580b6;
        mem[14'd1266] <= 32'h3b9f3f17;
        mem[14'd1267] <= 32'hbcbbfa80;
        mem[14'd1268] <= 32'hbcc5921d;
        mem[14'd1269] <= 32'h3ca3cc45;
        mem[14'd1270] <= 32'h3e63e900;
        mem[14'd1271] <= 32'h3e57a167;
        mem[14'd1272] <= 32'h3de14265;
        mem[14'd1273] <= 32'h3db74a61;
        mem[14'd1274] <= 32'h3e251bfb;
        mem[14'd1275] <= 32'h3dcbdca3;
        mem[14'd1276] <= 32'h3d7f8a40;
        mem[14'd1277] <= 32'hbea5f815;
        mem[14'd1278] <= 32'hbf1d0bc5;
        mem[14'd1279] <= 32'hbf3f3b9d;
        mem[14'd1280] <= 32'hbf133860;
        mem[14'd1281] <= 32'hbe60aab4;
        mem[14'd1282] <= 32'hbd0f9391;
        mem[14'd1283] <= 32'hbd9c506a;
        mem[14'd1284] <= 32'hbe2b5634;
        mem[14'd1285] <= 32'h3cd68e0b;
        mem[14'd1286] <= 32'h3e73585f;
        mem[14'd1287] <= 32'h3ecb8469;
        mem[14'd1288] <= 32'h3ea3ca8d;
        mem[14'd1289] <= 32'h3d284f38;
        mem[14'd1290] <= 32'hbb926bd8;
        mem[14'd1291] <= 32'hbc696013;
        mem[14'd1292] <= 32'h3c88bc33;
        mem[14'd1293] <= 32'h3a3bd503;
        mem[14'd1294] <= 32'hbb4443d5;
        mem[14'd1295] <= 32'hbcd1ba30;
        mem[14'd1296] <= 32'hbcf4cf02;
        mem[14'd1297] <= 32'h3e4e4037;
        mem[14'd1298] <= 32'h3e681978;
        mem[14'd1299] <= 32'h3e9ee7c0;
        mem[14'd1300] <= 32'h3e459050;
        mem[14'd1301] <= 32'h3e579a32;
        mem[14'd1302] <= 32'h3e19331c;
        mem[14'd1303] <= 32'h3e3a60d7;
        mem[14'd1304] <= 32'h3dadbc2b;
        mem[14'd1305] <= 32'hbe87b7c1;
        mem[14'd1306] <= 32'hbf2c07de;
        mem[14'd1307] <= 32'hbf314c10;
        mem[14'd1308] <= 32'hbf225c35;
        mem[14'd1309] <= 32'hbe2f648d;
        mem[14'd1310] <= 32'hbd7b7b90;
        mem[14'd1311] <= 32'hbe01109b;
        mem[14'd1312] <= 32'hbc4f30a5;
        mem[14'd1313] <= 32'h3e03667f;
        mem[14'd1314] <= 32'h3e256219;
        mem[14'd1315] <= 32'h3eb87f72;
        mem[14'd1316] <= 32'h3ea9ae0d;
        mem[14'd1317] <= 32'h3cebdfb9;
        mem[14'd1318] <= 32'hbc5e24d2;
        mem[14'd1319] <= 32'hbc72b868;
        mem[14'd1320] <= 32'h388dd9ca;
        mem[14'd1321] <= 32'h3a9eb102;
        mem[14'd1322] <= 32'h380082b3;
        mem[14'd1323] <= 32'hbd4430b3;
        mem[14'd1324] <= 32'h3ca9ef6d;
        mem[14'd1325] <= 32'h3e8684e7;
        mem[14'd1326] <= 32'h3defb213;
        mem[14'd1327] <= 32'h3e98bc58;
        mem[14'd1328] <= 32'h3e764e66;
        mem[14'd1329] <= 32'h3e77e2b9;
        mem[14'd1330] <= 32'h3e8028f3;
        mem[14'd1331] <= 32'h3da3b387;
        mem[14'd1332] <= 32'hbd8d3303;
        mem[14'd1333] <= 32'hbf0598ea;
        mem[14'd1334] <= 32'hbf435c44;
        mem[14'd1335] <= 32'hbf23a9b9;
        mem[14'd1336] <= 32'hbee033e9;
        mem[14'd1337] <= 32'hbe519f36;
        mem[14'd1338] <= 32'hbd4d9d74;
        mem[14'd1339] <= 32'hbd9832fa;
        mem[14'd1340] <= 32'h3e03b931;
        mem[14'd1341] <= 32'h3dd2ae89;
        mem[14'd1342] <= 32'h3e3cf40f;
        mem[14'd1343] <= 32'h3e999978;
        mem[14'd1344] <= 32'h3e6de06c;
        mem[14'd1345] <= 32'h3aa1c20a;
        mem[14'd1346] <= 32'hbc2c9e2b;
        mem[14'd1347] <= 32'h3bd170b5;
        mem[14'd1348] <= 32'h3ada98be;
        mem[14'd1349] <= 32'hbbba8733;
        mem[14'd1350] <= 32'hbbee78b9;
        mem[14'd1351] <= 32'hbd095b41;
        mem[14'd1352] <= 32'h3d1bb66b;
        mem[14'd1353] <= 32'h3e99be66;
        mem[14'd1354] <= 32'h3e5d5c14;
        mem[14'd1355] <= 32'h3e715b06;
        mem[14'd1356] <= 32'h3e898174;
        mem[14'd1357] <= 32'h3e877368;
        mem[14'd1358] <= 32'h3e8b70c5;
        mem[14'd1359] <= 32'h3dc36575;
        mem[14'd1360] <= 32'hbe87f44b;
        mem[14'd1361] <= 32'hbf2fc6ee;
        mem[14'd1362] <= 32'hbf2ecf87;
        mem[14'd1363] <= 32'hbee3bab0;
        mem[14'd1364] <= 32'hbe8006b6;
        mem[14'd1365] <= 32'hbd213424;
        mem[14'd1366] <= 32'h3c55faec;
        mem[14'd1367] <= 32'h3cfd0bcf;
        mem[14'd1368] <= 32'h3e3602be;
        mem[14'd1369] <= 32'h3e0534a9;
        mem[14'd1370] <= 32'h3e3c6efd;
        mem[14'd1371] <= 32'h3e52d1c5;
        mem[14'd1372] <= 32'h3daedd3e;
        mem[14'd1373] <= 32'hbd4c4e8d;
        mem[14'd1374] <= 32'hbd29f3fd;
        mem[14'd1375] <= 32'hbbef7b34;
        mem[14'd1376] <= 32'hbc8500c2;
        mem[14'd1377] <= 32'hbc07e0d8;
        mem[14'd1378] <= 32'h393b2844;
        mem[14'd1379] <= 32'hbd2a3a62;
        mem[14'd1380] <= 32'h3d64d0fb;
        mem[14'd1381] <= 32'h3e8090fd;
        mem[14'd1382] <= 32'h3e707c40;
        mem[14'd1383] <= 32'h3e3ff00f;
        mem[14'd1384] <= 32'h3e000f78;
        mem[14'd1385] <= 32'h3e86bff1;
        mem[14'd1386] <= 32'h3ebc3293;
        mem[14'd1387] <= 32'h3df5fa81;
        mem[14'd1388] <= 32'hbe5cc73b;
        mem[14'd1389] <= 32'hbf1cc600;
        mem[14'd1390] <= 32'hbf132a22;
        mem[14'd1391] <= 32'hbea3dde3;
        mem[14'd1392] <= 32'hbdb94d18;
        mem[14'd1393] <= 32'h3dbe94c3;
        mem[14'd1394] <= 32'h3c352265;
        mem[14'd1395] <= 32'h3d9d3ea3;
        mem[14'd1396] <= 32'h3dd7524c;
        mem[14'd1397] <= 32'h3d8aa19d;
        mem[14'd1398] <= 32'h3e2b68ea;
        mem[14'd1399] <= 32'h3dac0ddf;
        mem[14'd1400] <= 32'hbbab01fb;
        mem[14'd1401] <= 32'hbd34b011;
        mem[14'd1402] <= 32'hbc4f64c9;
        mem[14'd1403] <= 32'h3cb6e3ee;
        mem[14'd1404] <= 32'hbc20d082;
        mem[14'd1405] <= 32'hbbb49753;
        mem[14'd1406] <= 32'hbaf45483;
        mem[14'd1407] <= 32'hbd9ec2f1;
        mem[14'd1408] <= 32'hbcadc676;
        mem[14'd1409] <= 32'h3df65d8a;
        mem[14'd1410] <= 32'h3e2223e8;
        mem[14'd1411] <= 32'h3e19c3ad;
        mem[14'd1412] <= 32'h3e5d76be;
        mem[14'd1413] <= 32'h3e83e8cf;
        mem[14'd1414] <= 32'h3eb34a96;
        mem[14'd1415] <= 32'h3dd417dd;
        mem[14'd1416] <= 32'hbe876d27;
        mem[14'd1417] <= 32'hbf081f71;
        mem[14'd1418] <= 32'hbed5b727;
        mem[14'd1419] <= 32'hbe2e30d1;
        mem[14'd1420] <= 32'hbd63d432;
        mem[14'd1421] <= 32'hbc60dc80;
        mem[14'd1422] <= 32'hbc5aef7e;
        mem[14'd1423] <= 32'hb99bed5f;
        mem[14'd1424] <= 32'hbd16a19a;
        mem[14'd1425] <= 32'h3d880136;
        mem[14'd1426] <= 32'h3e30ae0b;
        mem[14'd1427] <= 32'h3d65c5d3;
        mem[14'd1428] <= 32'hbccb22b5;
        mem[14'd1429] <= 32'hbd1acf05;
        mem[14'd1430] <= 32'h3bd83f0e;
        mem[14'd1431] <= 32'h3bcf2b63;
        mem[14'd1432] <= 32'h39f5e118;
        mem[14'd1433] <= 32'hbbf3cc64;
        mem[14'd1434] <= 32'hbc520710;
        mem[14'd1435] <= 32'hbd6f82a2;
        mem[14'd1436] <= 32'hbd464736;
        mem[14'd1437] <= 32'h3ded3f77;
        mem[14'd1438] <= 32'h3e4555d9;
        mem[14'd1439] <= 32'h3e57b086;
        mem[14'd1440] <= 32'h3e59f5b3;
        mem[14'd1441] <= 32'h3e25a41f;
        mem[14'd1442] <= 32'h3e973332;
        mem[14'd1443] <= 32'h3e93a74c;
        mem[14'd1444] <= 32'h3e0cc26f;
        mem[14'd1445] <= 32'hbe1498d4;
        mem[14'd1446] <= 32'hbe5e2989;
        mem[14'd1447] <= 32'hbe0aece6;
        mem[14'd1448] <= 32'hbdc13512;
        mem[14'd1449] <= 32'h3cbf1778;
        mem[14'd1450] <= 32'hbc81547b;
        mem[14'd1451] <= 32'hbd783e92;
        mem[14'd1452] <= 32'h3c608d36;
        mem[14'd1453] <= 32'h3dadda06;
        mem[14'd1454] <= 32'h3e0e813a;
        mem[14'd1455] <= 32'h3caa0f5c;
        mem[14'd1456] <= 32'hbd0fc990;
        mem[14'd1457] <= 32'hbbdcf089;
        mem[14'd1458] <= 32'h3b700bf3;
        mem[14'd1459] <= 32'hbc8bb32d;
        mem[14'd1460] <= 32'h3c4d0a8a;
        mem[14'd1461] <= 32'hbb60a5e8;
        mem[14'd1462] <= 32'h3c8cbe02;
        mem[14'd1463] <= 32'hbd0ed88e;
        mem[14'd1464] <= 32'hbc5c0971;
        mem[14'd1465] <= 32'h3e19d22e;
        mem[14'd1466] <= 32'h3e1bbc9e;
        mem[14'd1467] <= 32'h3e02b96d;
        mem[14'd1468] <= 32'h3e14ab9c;
        mem[14'd1469] <= 32'h3e26e83e;
        mem[14'd1470] <= 32'h3eae61b7;
        mem[14'd1471] <= 32'h3ed3c5b3;
        mem[14'd1472] <= 32'h3eb527e3;
        mem[14'd1473] <= 32'h3e0f295e;
        mem[14'd1474] <= 32'hbcf8eb16;
        mem[14'd1475] <= 32'hbba120c6;
        mem[14'd1476] <= 32'hbd6e5fb9;
        mem[14'd1477] <= 32'hbcd6b9bb;
        mem[14'd1478] <= 32'hbe02bc27;
        mem[14'd1479] <= 32'hbe0afff6;
        mem[14'd1480] <= 32'hbdb7fe72;
        mem[14'd1481] <= 32'h3d4de9d3;
        mem[14'd1482] <= 32'h3d68b485;
        mem[14'd1483] <= 32'hbd8c68d2;
        mem[14'd1484] <= 32'hbd80df83;
        mem[14'd1485] <= 32'hbcc139c9;
        mem[14'd1486] <= 32'h3c0fd97c;
        mem[14'd1487] <= 32'hbc44e5bb;
        mem[14'd1488] <= 32'hbc491666;
        mem[14'd1489] <= 32'hbb4b5f20;
        mem[14'd1490] <= 32'hbc0a9d2f;
        mem[14'd1491] <= 32'hbd3ee1e2;
        mem[14'd1492] <= 32'hbd5a77ca;
        mem[14'd1493] <= 32'h3d9bc361;
        mem[14'd1494] <= 32'h3e079951;
        mem[14'd1495] <= 32'h3de6c82e;
        mem[14'd1496] <= 32'h3d07ede0;
        mem[14'd1497] <= 32'h3d6d1f09;
        mem[14'd1498] <= 32'h3e56faee;
        mem[14'd1499] <= 32'h3ea7d288;
        mem[14'd1500] <= 32'h3e86f769;
        mem[14'd1501] <= 32'h3da04d4d;
        mem[14'd1502] <= 32'h3c415579;
        mem[14'd1503] <= 32'h3c15c829;
        mem[14'd1504] <= 32'hbb0acc51;
        mem[14'd1505] <= 32'hbe2354f2;
        mem[14'd1506] <= 32'hbe2471c0;
        mem[14'd1507] <= 32'hbe3d4388;
        mem[14'd1508] <= 32'hbd8b2532;
        mem[14'd1509] <= 32'h3bafb737;
        mem[14'd1510] <= 32'hbc7a709b;
        mem[14'd1511] <= 32'hbd69736e;
        mem[14'd1512] <= 32'hbd55a48e;
        mem[14'd1513] <= 32'hbc0e81e7;
        mem[14'd1514] <= 32'h3ad208e6;
        mem[14'd1515] <= 32'hbc12ac58;
        mem[14'd1516] <= 32'hbc07c06a;
        mem[14'd1517] <= 32'h3b15f571;
        mem[14'd1518] <= 32'h3c69b65b;
        mem[14'd1519] <= 32'hbc4839fc;
        mem[14'd1520] <= 32'hbe270b26;
        mem[14'd1521] <= 32'hbc97018f;
        mem[14'd1522] <= 32'h3d866fc5;
        mem[14'd1523] <= 32'h3d9a568a;
        mem[14'd1524] <= 32'h3e1ee00c;
        mem[14'd1525] <= 32'h3e11a3a1;
        mem[14'd1526] <= 32'h3e18e9f6;
        mem[14'd1527] <= 32'h3e3972af;
        mem[14'd1528] <= 32'h3e48f946;
        mem[14'd1529] <= 32'h3eadd611;
        mem[14'd1530] <= 32'h3e290792;
        mem[14'd1531] <= 32'h3dfb3440;
        mem[14'd1532] <= 32'h3d1145ea;
        mem[14'd1533] <= 32'hbc8a9176;
        mem[14'd1534] <= 32'hbdccd9cf;
        mem[14'd1535] <= 32'hbde6353d;
        mem[14'd1536] <= 32'hbdefd216;
        mem[14'd1537] <= 32'hbdc5ab20;
        mem[14'd1538] <= 32'hbcabb8a4;
        mem[14'd1539] <= 32'hbd277ae8;
        mem[14'd1540] <= 32'hbd10e15c;
        mem[14'd1541] <= 32'hbb77fb4d;
        mem[14'd1542] <= 32'hbb57fc1f;
        mem[14'd1543] <= 32'h3b1127af;
        mem[14'd1544] <= 32'hb91c5ec9;
        mem[14'd1545] <= 32'hbc0938e9;
        mem[14'd1546] <= 32'h3b90c5fc;
        mem[14'd1547] <= 32'hbd0c5304;
        mem[14'd1548] <= 32'hbdf3c671;
        mem[14'd1549] <= 32'hbdce0ebc;
        mem[14'd1550] <= 32'hbc7bfae8;
        mem[14'd1551] <= 32'h3d4e5ce2;
        mem[14'd1552] <= 32'h3db34965;
        mem[14'd1553] <= 32'h3e674d98;
        mem[14'd1554] <= 32'h3ea99bbc;
        mem[14'd1555] <= 32'h3ead7779;
        mem[14'd1556] <= 32'h3e9bd74f;
        mem[14'd1557] <= 32'h3e9ad443;
        mem[14'd1558] <= 32'h3e7d12c2;
        mem[14'd1559] <= 32'h3e143ecb;
        mem[14'd1560] <= 32'h3ce4fbad;
        mem[14'd1561] <= 32'hba4807b2;
        mem[14'd1562] <= 32'hbe3af1de;
        mem[14'd1563] <= 32'hbe7e303c;
        mem[14'd1564] <= 32'hbe65a02d;
        mem[14'd1565] <= 32'hbe09649e;
        mem[14'd1566] <= 32'hbd462a17;
        mem[14'd1567] <= 32'hbce5cc6e;
        mem[14'd1568] <= 32'hbd166510;
        mem[14'd1569] <= 32'h3c713b81;
        mem[14'd1570] <= 32'hbb005c32;
        mem[14'd1571] <= 32'h3bf29e13;
        mem[14'd1572] <= 32'hb93232c8;
        mem[14'd1573] <= 32'hbb3e65f9;
        mem[14'd1574] <= 32'hbb6a0add;
        mem[14'd1575] <= 32'h3be3bc06;
        mem[14'd1576] <= 32'hbca65864;
        mem[14'd1577] <= 32'hbd39b799;
        mem[14'd1578] <= 32'hbdbc5946;
        mem[14'd1579] <= 32'hbdcf405f;
        mem[14'd1580] <= 32'hbdde8e6c;
        mem[14'd1581] <= 32'hbd37bc9e;
        mem[14'd1582] <= 32'hbd0979e9;
        mem[14'd1583] <= 32'h3c7d717f;
        mem[14'd1584] <= 32'h3e10da1f;
        mem[14'd1585] <= 32'h3e0ac291;
        mem[14'd1586] <= 32'h3d8f9b0e;
        mem[14'd1587] <= 32'hbcb34bcd;
        mem[14'd1588] <= 32'hbdd099e8;
        mem[14'd1589] <= 32'hbe1db2f3;
        mem[14'd1590] <= 32'hbe558b22;
        mem[14'd1591] <= 32'hbe58e5dd;
        mem[14'd1592] <= 32'hbe3e8e28;
        mem[14'd1593] <= 32'hbddb5940;
        mem[14'd1594] <= 32'hbd838c2b;
        mem[14'd1595] <= 32'hbaed9dc7;
        mem[14'd1596] <= 32'h3b8bd1cc;
        mem[14'd1597] <= 32'h3bd2ce2e;
        mem[14'd1598] <= 32'hbba6df4d;
        mem[14'd1599] <= 32'hbc62ed62;
        mem[14'd1600] <= 32'h3b884204;
        mem[14'd1601] <= 32'h3ca72879;
        mem[14'd1602] <= 32'hba838e10;
        mem[14'd1603] <= 32'h3be2207b;
        mem[14'd1604] <= 32'h3b8eeb1a;
        mem[14'd1605] <= 32'hbc756868;
        mem[14'd1606] <= 32'hbd5da64a;
        mem[14'd1607] <= 32'hbda3c9ef;
        mem[14'd1608] <= 32'hbe07e4fd;
        mem[14'd1609] <= 32'hbe5774e9;
        mem[14'd1610] <= 32'hbe861be4;
        mem[14'd1611] <= 32'hbe82d710;
        mem[14'd1612] <= 32'hbe96fa40;
        mem[14'd1613] <= 32'hbe82afaf;
        mem[14'd1614] <= 32'hbe93b1d2;
        mem[14'd1615] <= 32'hbe73ddcf;
        mem[14'd1616] <= 32'hbe47f852;
        mem[14'd1617] <= 32'hbe2edaac;
        mem[14'd1618] <= 32'hbe207c0a;
        mem[14'd1619] <= 32'hbdcf429d;
        mem[14'd1620] <= 32'hbdbe5b61;
        mem[14'd1621] <= 32'hbdb29b9d;
        mem[14'd1622] <= 32'hbcf218c2;
        mem[14'd1623] <= 32'hb9a7b0f3;
        mem[14'd1624] <= 32'hbc0d7d12;
        mem[14'd1625] <= 32'h3c11c84a;
        mem[14'd1626] <= 32'hbc2ec96e;
        mem[14'd1627] <= 32'h3bf3cf8f;
        mem[14'd1628] <= 32'h3c578b79;
        mem[14'd1629] <= 32'h3b3d20af;
        mem[14'd1630] <= 32'hbbf6316e;
        mem[14'd1631] <= 32'hbc86dd4e;
        mem[14'd1632] <= 32'h3c121d42;
        mem[14'd1633] <= 32'hbc7c68d4;
        mem[14'd1634] <= 32'hba993b6c;
        mem[14'd1635] <= 32'hbd158a9b;
        mem[14'd1636] <= 32'hbccf1f44;
        mem[14'd1637] <= 32'hbd961499;
        mem[14'd1638] <= 32'hbd96c68a;
        mem[14'd1639] <= 32'hbcf55a7e;
        mem[14'd1640] <= 32'hbcf05643;
        mem[14'd1641] <= 32'hbd7caca8;
        mem[14'd1642] <= 32'hbda08523;
        mem[14'd1643] <= 32'hbd7a9db5;
        mem[14'd1644] <= 32'hbd4a713d;
        mem[14'd1645] <= 32'hbd43145b;
        mem[14'd1646] <= 32'hbd1f7ade;
        mem[14'd1647] <= 32'hbbfca355;
        mem[14'd1648] <= 32'hbd0f8255;
        mem[14'd1649] <= 32'hbd0f785b;
        mem[14'd1650] <= 32'hbc5c8693;
        mem[14'd1651] <= 32'hbc02e93c;
        mem[14'd1652] <= 32'h38652b37;
        mem[14'd1653] <= 32'h3cab0563;
        mem[14'd1654] <= 32'h399baa17;
        mem[14'd1655] <= 32'h3aa13e21;
        mem[14'd1656] <= 32'hbc1738f0;
        mem[14'd1657] <= 32'h3c1ed8db;
        mem[14'd1658] <= 32'hbb90f1ad;
        mem[14'd1659] <= 32'hbb2c064f;
        mem[14'd1660] <= 32'hbbef8e86;
        mem[14'd1661] <= 32'hbc9daa43;
        mem[14'd1662] <= 32'hbb981ba1;
        mem[14'd1663] <= 32'h390786e8;
        mem[14'd1664] <= 32'h3c330e2a;
        mem[14'd1665] <= 32'h3a35349b;
        mem[14'd1666] <= 32'h3c5e6dfb;
        mem[14'd1667] <= 32'hbc5d2f07;
        mem[14'd1668] <= 32'hbc83cb24;
        mem[14'd1669] <= 32'hbc324909;
        mem[14'd1670] <= 32'hbc821ad2;
        mem[14'd1671] <= 32'hbc4ed198;
        mem[14'd1672] <= 32'hbc936957;
        mem[14'd1673] <= 32'hbc57e707;
        mem[14'd1674] <= 32'hbc341d20;
        mem[14'd1675] <= 32'hbc9df94b;
        mem[14'd1676] <= 32'hbba99e2b;
        mem[14'd1677] <= 32'hb9efbed0;
        mem[14'd1678] <= 32'hbca5d7e9;
        mem[14'd1679] <= 32'hbb51f03e;
        mem[14'd1680] <= 32'hbc68fb3b;
        mem[14'd1681] <= 32'h3ca771eb;
        mem[14'd1682] <= 32'hbc204975;
        mem[14'd1683] <= 32'h3c52a493;
        mem[14'd1684] <= 32'hbb1a7634;
        mem[14'd1685] <= 32'hbb7ccb09;
        mem[14'd1686] <= 32'hba184779;
        mem[14'd1687] <= 32'hbb198344;
        mem[14'd1688] <= 32'h3abc2f4a;
        mem[14'd1689] <= 32'hbc483147;
        mem[14'd1690] <= 32'h3b3b9ddc;
        mem[14'd1691] <= 32'hbc062b66;
        mem[14'd1692] <= 32'h3c2eb3fc;
        mem[14'd1693] <= 32'hbb6054be;
        mem[14'd1694] <= 32'h391943d1;
        mem[14'd1695] <= 32'hbbee09ce;
        mem[14'd1696] <= 32'h3bddc371;
        mem[14'd1697] <= 32'hbba6b41d;
        mem[14'd1698] <= 32'h3b7a5197;
        mem[14'd1699] <= 32'h3b37b94f;
        mem[14'd1700] <= 32'h3b194316;
        mem[14'd1701] <= 32'h3c881a8b;
        mem[14'd1702] <= 32'hbbd85707;
        mem[14'd1703] <= 32'hbb5fba41;
        mem[14'd1704] <= 32'h3b72eb63;
        mem[14'd1705] <= 32'hbc406e0e;
        mem[14'd1706] <= 32'h3c968fdf;
        mem[14'd1707] <= 32'h3be43b6f;
        mem[14'd1708] <= 32'hbc2f1006;
        mem[14'd1709] <= 32'h3b74e603;
        mem[14'd1710] <= 32'hbc2406f9;
        mem[14'd1711] <= 32'hbcae0baf;
        mem[14'd1712] <= 32'hbc7dece7;
        mem[14'd1713] <= 32'h3b15a39c;
        mem[14'd1714] <= 32'h3b017d7f;
        mem[14'd1715] <= 32'hbc0f8017;
        mem[14'd1716] <= 32'h3c5f709b;
        mem[14'd1717] <= 32'hbb56fe92;
        mem[14'd1718] <= 32'h3bdcb1fd;
        mem[14'd1719] <= 32'hbc837594;
        mem[14'd1720] <= 32'h3b28ee79;
        mem[14'd1721] <= 32'hbc97737e;
        mem[14'd1722] <= 32'h3c1e431b;
        mem[14'd1723] <= 32'hbbc61509;
        mem[14'd1724] <= 32'h3c21167b;
        mem[14'd1725] <= 32'hbc73606b;
        mem[14'd1726] <= 32'h3cc33408;
        mem[14'd1727] <= 32'h3d06cac8;
        mem[14'd1728] <= 32'h3c2c8463;
        mem[14'd1729] <= 32'h3bf78254;
        mem[14'd1730] <= 32'hbc408142;
        mem[14'd1731] <= 32'hbc9ae351;
        mem[14'd1732] <= 32'hbb49e858;
        mem[14'd1733] <= 32'hbb68b55f;
        mem[14'd1734] <= 32'h3c0f4449;
        mem[14'd1735] <= 32'h3bd40996;
        mem[14'd1736] <= 32'hbb85ea55;
        mem[14'd1737] <= 32'h3ac03ff5;
        mem[14'd1738] <= 32'h3c8fba07;
        mem[14'd1739] <= 32'h3bc5ff59;
        mem[14'd1740] <= 32'hbbadfca2;
        mem[14'd1741] <= 32'hbc0d21bf;
        mem[14'd1742] <= 32'h3ad90ea6;
        mem[14'd1743] <= 32'h3bcf8a65;
        mem[14'd1744] <= 32'hbb74673e;
        mem[14'd1745] <= 32'h3c45c3b9;
        mem[14'd1746] <= 32'h3c238f2a;
        mem[14'd1747] <= 32'hbb913638;
        mem[14'd1748] <= 32'hbca7728f;
        mem[14'd1749] <= 32'hbcc302bb;
        mem[14'd1750] <= 32'hbc82f379;
        mem[14'd1751] <= 32'hbd06b825;
        mem[14'd1752] <= 32'h3b135855;
        mem[14'd1753] <= 32'h3d406499;
        mem[14'd1754] <= 32'h3d68cf5a;
        mem[14'd1755] <= 32'h3df4ed3c;
        mem[14'd1756] <= 32'h3da5f62b;
        mem[14'd1757] <= 32'h3d17b00b;
        mem[14'd1758] <= 32'hbc8b880e;
        mem[14'd1759] <= 32'h3a9ad679;
        mem[14'd1760] <= 32'hbbbf287c;
        mem[14'd1761] <= 32'hbac89b2b;
        mem[14'd1762] <= 32'h3c4624fc;
        mem[14'd1763] <= 32'hbc5cd821;
        mem[14'd1764] <= 32'hbc8d185f;
        mem[14'd1765] <= 32'hbb4d7c8b;
        mem[14'd1766] <= 32'h39cd35c6;
        mem[14'd1767] <= 32'hbc0b1a3d;
        mem[14'd1768] <= 32'h3bb23c29;
        mem[14'd1769] <= 32'h3adadb78;
        mem[14'd1770] <= 32'h3b2ccb6f;
        mem[14'd1771] <= 32'h3c6e5ad9;
        mem[14'd1772] <= 32'hba5fd5c3;
        mem[14'd1773] <= 32'hbbaa765d;
        mem[14'd1774] <= 32'hbc9242f2;
        mem[14'd1775] <= 32'hbcf3113b;
        mem[14'd1776] <= 32'hbd326cd4;
        mem[14'd1777] <= 32'hbd997aad;
        mem[14'd1778] <= 32'hbdc8b323;
        mem[14'd1779] <= 32'hbe2970a6;
        mem[14'd1780] <= 32'hbd9dd17d;
        mem[14'd1781] <= 32'hbce34454;
        mem[14'd1782] <= 32'hbd0ff9de;
        mem[14'd1783] <= 32'h3d6007a7;
        mem[14'd1784] <= 32'h3d6f12f6;
        mem[14'd1785] <= 32'hbd3faddf;
        mem[14'd1786] <= 32'hbde9877a;
        mem[14'd1787] <= 32'hbd8083e6;
        mem[14'd1788] <= 32'hbd84853c;
        mem[14'd1789] <= 32'hbd855ad9;
        mem[14'd1790] <= 32'hbd726dd6;
        mem[14'd1791] <= 32'hbccf37bf;
        mem[14'd1792] <= 32'hbcbe838d;
        mem[14'd1793] <= 32'hbbf51909;
        mem[14'd1794] <= 32'hbcbe4e90;
        mem[14'd1795] <= 32'h3b8e1d45;
        mem[14'd1796] <= 32'hbbedd51e;
        mem[14'd1797] <= 32'h3b1a790b;
        mem[14'd1798] <= 32'h3b8f3a0d;
        mem[14'd1799] <= 32'h3c5bbacf;
        mem[14'd1800] <= 32'hbc588059;
        mem[14'd1801] <= 32'h3b1c8be3;
        mem[14'd1802] <= 32'hbc70514d;
        mem[14'd1803] <= 32'hbd1a1862;
        mem[14'd1804] <= 32'hbcc496e8;
        mem[14'd1805] <= 32'hbdbcd88a;
        mem[14'd1806] <= 32'hbd9f0559;
        mem[14'd1807] <= 32'hbe18b975;
        mem[14'd1808] <= 32'hbd0a7f0f;
        mem[14'd1809] <= 32'h3e0a54c8;
        mem[14'd1810] <= 32'h3e1023ec;
        mem[14'd1811] <= 32'h3e008232;
        mem[14'd1812] <= 32'h3d7ecac8;
        mem[14'd1813] <= 32'hbd5182b5;
        mem[14'd1814] <= 32'hbd2b532d;
        mem[14'd1815] <= 32'h3daa55a2;
        mem[14'd1816] <= 32'h3dbed573;
        mem[14'd1817] <= 32'h3da71af4;
        mem[14'd1818] <= 32'h3cc83b62;
        mem[14'd1819] <= 32'h3c23965b;
        mem[14'd1820] <= 32'hbda5cd98;
        mem[14'd1821] <= 32'hbd238f2e;
        mem[14'd1822] <= 32'h3be721ec;
        mem[14'd1823] <= 32'hbc19f58f;
        mem[14'd1824] <= 32'hbbbafdf8;
        mem[14'd1825] <= 32'hbaa2c0be;
        mem[14'd1826] <= 32'hbba17558;
        mem[14'd1827] <= 32'h3c43334e;
        mem[14'd1828] <= 32'h3c56cf85;
        mem[14'd1829] <= 32'h3d3bb9e0;
        mem[14'd1830] <= 32'hbb8c1b79;
        mem[14'd1831] <= 32'hbd3f676e;
        mem[14'd1832] <= 32'hbe344bdd;
        mem[14'd1833] <= 32'hbe513f7f;
        mem[14'd1834] <= 32'hbe398be4;
        mem[14'd1835] <= 32'hbe409c16;
        mem[14'd1836] <= 32'hbdb6717b;
        mem[14'd1837] <= 32'h3cfa2e58;
        mem[14'd1838] <= 32'h3db4d344;
        mem[14'd1839] <= 32'h3e1c07a3;
        mem[14'd1840] <= 32'hbcbf1606;
        mem[14'd1841] <= 32'hbe0c394e;
        mem[14'd1842] <= 32'hbbb9e876;
        mem[14'd1843] <= 32'h3d7d827e;
        mem[14'd1844] <= 32'h3df09193;
        mem[14'd1845] <= 32'h3e65c177;
        mem[14'd1846] <= 32'h3e50646b;
        mem[14'd1847] <= 32'h3dfb2377;
        mem[14'd1848] <= 32'hb986fcee;
        mem[14'd1849] <= 32'hbd645242;
        mem[14'd1850] <= 32'hbc9d42a6;
        mem[14'd1851] <= 32'hbc19bf32;
        mem[14'd1852] <= 32'hbb96615c;
        mem[14'd1853] <= 32'h3b08870a;
        mem[14'd1854] <= 32'h3b12e14f;
        mem[14'd1855] <= 32'h3c071a93;
        mem[14'd1856] <= 32'h3b93d57d;
        mem[14'd1857] <= 32'hbc662522;
        mem[14'd1858] <= 32'hbd2b13df;
        mem[14'd1859] <= 32'hbe16351f;
        mem[14'd1860] <= 32'hbe7cc3dc;
        mem[14'd1861] <= 32'hbe8b3001;
        mem[14'd1862] <= 32'hbe4f68e3;
        mem[14'd1863] <= 32'hbde8419b;
        mem[14'd1864] <= 32'hbe327783;
        mem[14'd1865] <= 32'hbe1b980e;
        mem[14'd1866] <= 32'hbe1331b2;
        mem[14'd1867] <= 32'hbe5cf418;
        mem[14'd1868] <= 32'hbe6c7ab6;
        mem[14'd1869] <= 32'hbe834b78;
        mem[14'd1870] <= 32'hbdc31802;
        mem[14'd1871] <= 32'hbd9ebdf1;
        mem[14'd1872] <= 32'h3d8482f9;
        mem[14'd1873] <= 32'h3db8f152;
        mem[14'd1874] <= 32'h3db4bbd8;
        mem[14'd1875] <= 32'h3d1fb96e;
        mem[14'd1876] <= 32'hbd2b326d;
        mem[14'd1877] <= 32'hbd73d9cf;
        mem[14'd1878] <= 32'hbc6bc123;
        mem[14'd1879] <= 32'hbc8fcced;
        mem[14'd1880] <= 32'hbc3d536d;
        mem[14'd1881] <= 32'hbc8631e0;
        mem[14'd1882] <= 32'h3b9d70a8;
        mem[14'd1883] <= 32'hbc269f5f;
        mem[14'd1884] <= 32'hbc27b55b;
        mem[14'd1885] <= 32'hbd93ed9c;
        mem[14'd1886] <= 32'hbe2cbb05;
        mem[14'd1887] <= 32'hbe2cf22e;
        mem[14'd1888] <= 32'hbe9a4bb7;
        mem[14'd1889] <= 32'hbe919878;
        mem[14'd1890] <= 32'hbe6eaf6f;
        mem[14'd1891] <= 32'hbe576c2a;
        mem[14'd1892] <= 32'hbdd5f5b1;
        mem[14'd1893] <= 32'hbe25612b;
        mem[14'd1894] <= 32'hbe06dcc9;
        mem[14'd1895] <= 32'hbe9bfc64;
        mem[14'd1896] <= 32'hbe693b51;
        mem[14'd1897] <= 32'hbe55c21d;
        mem[14'd1898] <= 32'hbe33c1d9;
        mem[14'd1899] <= 32'hbd405674;
        mem[14'd1900] <= 32'h3d57a548;
        mem[14'd1901] <= 32'hbc9bb640;
        mem[14'd1902] <= 32'hbc313363;
        mem[14'd1903] <= 32'hbdd7b97f;
        mem[14'd1904] <= 32'hbe45b93a;
        mem[14'd1905] <= 32'hbdd6c1a5;
        mem[14'd1906] <= 32'hbbf72d32;
        mem[14'd1907] <= 32'hbbef0b30;
        mem[14'd1908] <= 32'hbb805d38;
        mem[14'd1909] <= 32'hbc650627;
        mem[14'd1910] <= 32'hbbc08a9f;
        mem[14'd1911] <= 32'hbc2075e6;
        mem[14'd1912] <= 32'hbd01ddff;
        mem[14'd1913] <= 32'hbdb3caa0;
        mem[14'd1914] <= 32'hbe148ea5;
        mem[14'd1915] <= 32'hbe3b08eb;
        mem[14'd1916] <= 32'hbe97e56e;
        mem[14'd1917] <= 32'hbea70438;
        mem[14'd1918] <= 32'hbe88734d;
        mem[14'd1919] <= 32'hbe48f4ee;
        mem[14'd1920] <= 32'hbd82e6b7;
        mem[14'd1921] <= 32'hbc6ab5b5;
        mem[14'd1922] <= 32'hbc8b1687;
        mem[14'd1923] <= 32'h3c39e45d;
        mem[14'd1924] <= 32'hbe20884d;
        mem[14'd1925] <= 32'h3cec7a27;
        mem[14'd1926] <= 32'hbdac062d;
        mem[14'd1927] <= 32'hbdcc7b8c;
        mem[14'd1928] <= 32'hbe1f9395;
        mem[14'd1929] <= 32'hbe39bf48;
        mem[14'd1930] <= 32'hbe47fe2d;
        mem[14'd1931] <= 32'hbea04b66;
        mem[14'd1932] <= 32'hbe9365a2;
        mem[14'd1933] <= 32'hbde08aa4;
        mem[14'd1934] <= 32'hbc5cb18b;
        mem[14'd1935] <= 32'h3b5f1280;
        mem[14'd1936] <= 32'hbc0b8e07;
        mem[14'd1937] <= 32'h3c31c8f6;
        mem[14'd1938] <= 32'hbc382b77;
        mem[14'd1939] <= 32'hbb5abf57;
        mem[14'd1940] <= 32'hbd509c49;
        mem[14'd1941] <= 32'hbe1264b0;
        mem[14'd1942] <= 32'hbe1b754b;
        mem[14'd1943] <= 32'hbe16d73f;
        mem[14'd1944] <= 32'hbe68807a;
        mem[14'd1945] <= 32'hbe868daf;
        mem[14'd1946] <= 32'hbe3027a8;
        mem[14'd1947] <= 32'hbd3d083a;
        mem[14'd1948] <= 32'hbd600b20;
        mem[14'd1949] <= 32'h3d260e77;
        mem[14'd1950] <= 32'h3e47fcd0;
        mem[14'd1951] <= 32'h3ecc7646;
        mem[14'd1952] <= 32'h3dff9092;
        mem[14'd1953] <= 32'h399b1c69;
        mem[14'd1954] <= 32'hbdf968aa;
        mem[14'd1955] <= 32'hbe6cd45a;
        mem[14'd1956] <= 32'hbe929c6b;
        mem[14'd1957] <= 32'hbe9083f6;
        mem[14'd1958] <= 32'hbea504d0;
        mem[14'd1959] <= 32'hbeabd88d;
        mem[14'd1960] <= 32'hbe5c53c8;
        mem[14'd1961] <= 32'hbdaecece;
        mem[14'd1962] <= 32'hbc35482a;
        mem[14'd1963] <= 32'hbbd3b9c8;
        mem[14'd1964] <= 32'hbc0cef5a;
        mem[14'd1965] <= 32'hbbb46748;
        mem[14'd1966] <= 32'hbc596b34;
        mem[14'd1967] <= 32'hbca6e0c8;
        mem[14'd1968] <= 32'hbd46780a;
        mem[14'd1969] <= 32'hbe01f980;
        mem[14'd1970] <= 32'hbe3ab3cd;
        mem[14'd1971] <= 32'hbe3e55a3;
        mem[14'd1972] <= 32'hbe35e277;
        mem[14'd1973] <= 32'hbe570e4f;
        mem[14'd1974] <= 32'hbd8c8f7e;
        mem[14'd1975] <= 32'hbb8871e3;
        mem[14'd1976] <= 32'hb9b37265;
        mem[14'd1977] <= 32'h3e52a075;
        mem[14'd1978] <= 32'h3f0479f3;
        mem[14'd1979] <= 32'h3f2af5d1;
        mem[14'd1980] <= 32'h3e8729dc;
        mem[14'd1981] <= 32'h3d2825b6;
        mem[14'd1982] <= 32'hbe3998ed;
        mem[14'd1983] <= 32'hbe5da5c3;
        mem[14'd1984] <= 32'hbea912bd;
        mem[14'd1985] <= 32'hbe98bb29;
        mem[14'd1986] <= 32'hbe9370bf;
        mem[14'd1987] <= 32'hbe8594e2;
        mem[14'd1988] <= 32'hbe404df8;
        mem[14'd1989] <= 32'hbd79a182;
        mem[14'd1990] <= 32'hbc81ea95;
        mem[14'd1991] <= 32'hbc41a6aa;
        mem[14'd1992] <= 32'h3bad9090;
        mem[14'd1993] <= 32'hbc40ada5;
        mem[14'd1994] <= 32'hbbce4d1d;
        mem[14'd1995] <= 32'hbd005d53;
        mem[14'd1996] <= 32'hbcbcfd12;
        mem[14'd1997] <= 32'hbda9be14;
        mem[14'd1998] <= 32'hbe1f1f11;
        mem[14'd1999] <= 32'hbe20a022;
        mem[14'd2000] <= 32'hbe404884;
        mem[14'd2001] <= 32'hbe4aeb5d;
        mem[14'd2002] <= 32'hbe1f91b0;
        mem[14'd2003] <= 32'hbe15efd5;
        mem[14'd2004] <= 32'hbd80fe67;
        mem[14'd2005] <= 32'h3e89b892;
        mem[14'd2006] <= 32'h3f2d7a41;
        mem[14'd2007] <= 32'h3f2c0b6f;
        mem[14'd2008] <= 32'h3e489966;
        mem[14'd2009] <= 32'hbd3ffe63;
        mem[14'd2010] <= 32'hbd2e81f9;
        mem[14'd2011] <= 32'hbe2bc141;
        mem[14'd2012] <= 32'hbe5bea1d;
        mem[14'd2013] <= 32'hbe4de130;
        mem[14'd2014] <= 32'hbe1365d3;
        mem[14'd2015] <= 32'hbdfc00ae;
        mem[14'd2016] <= 32'hbd9bf6d0;
        mem[14'd2017] <= 32'hbd068cf4;
        mem[14'd2018] <= 32'h3a9adc8a;
        mem[14'd2019] <= 32'h3c86b092;
        mem[14'd2020] <= 32'h3cbb5395;
        mem[14'd2021] <= 32'hba5b9988;
        mem[14'd2022] <= 32'h3be04f0a;
        mem[14'd2023] <= 32'hbbbb6c4c;
        mem[14'd2024] <= 32'h3c01ff49;
        mem[14'd2025] <= 32'hbd2942d3;
        mem[14'd2026] <= 32'hbd6ac0c8;
        mem[14'd2027] <= 32'hbd80437c;
        mem[14'd2028] <= 32'hbdd8a980;
        mem[14'd2029] <= 32'hbe15291e;
        mem[14'd2030] <= 32'hbe992725;
        mem[14'd2031] <= 32'hbece1ba6;
        mem[14'd2032] <= 32'hbd9ff5f9;
        mem[14'd2033] <= 32'h3e9068dd;
        mem[14'd2034] <= 32'h3f50cff0;
        mem[14'd2035] <= 32'h3f014053;
        mem[14'd2036] <= 32'h3dd4ba87;
        mem[14'd2037] <= 32'h3d95bdf3;
        mem[14'd2038] <= 32'hbcc6a267;
        mem[14'd2039] <= 32'hbe38d0fb;
        mem[14'd2040] <= 32'hbe2acd19;
        mem[14'd2041] <= 32'hbdcd41f3;
        mem[14'd2042] <= 32'hbdb21607;
        mem[14'd2043] <= 32'hbd48f71c;
        mem[14'd2044] <= 32'hbd1d5e98;
        mem[14'd2045] <= 32'hbc57b1b7;
        mem[14'd2046] <= 32'h3b61283b;
        mem[14'd2047] <= 32'h3c49724a;
        mem[14'd2048] <= 32'h3c774272;
        mem[14'd2049] <= 32'hbc4187bc;
        mem[14'd2050] <= 32'h3bbd7cd0;
        mem[14'd2051] <= 32'hba88f2eb;
        mem[14'd2052] <= 32'h3c753013;
        mem[14'd2053] <= 32'hbd453b70;
        mem[14'd2054] <= 32'hbd41424f;
        mem[14'd2055] <= 32'hbd9d595c;
        mem[14'd2056] <= 32'hbd3a0a87;
        mem[14'd2057] <= 32'hbe3bef55;
        mem[14'd2058] <= 32'hbf051ad6;
        mem[14'd2059] <= 32'hbf10ce8a;
        mem[14'd2060] <= 32'hbddbd89b;
        mem[14'd2061] <= 32'h3ea0b5ed;
        mem[14'd2062] <= 32'h3f1fb1e1;
        mem[14'd2063] <= 32'h3ec76af9;
        mem[14'd2064] <= 32'h3e17e66a;
        mem[14'd2065] <= 32'h3dee494d;
        mem[14'd2066] <= 32'hbe6b7e24;
        mem[14'd2067] <= 32'hbe804429;
        mem[14'd2068] <= 32'hbe3b5af8;
        mem[14'd2069] <= 32'hbdd51f40;
        mem[14'd2070] <= 32'hbdba8c1b;
        mem[14'd2071] <= 32'hbd9cd616;
        mem[14'd2072] <= 32'hbd7903f0;
        mem[14'd2073] <= 32'hbd32f7d5;
        mem[14'd2074] <= 32'hbccfe5e7;
        mem[14'd2075] <= 32'hbb910594;
        mem[14'd2076] <= 32'h3ba18957;
        mem[14'd2077] <= 32'hbc395220;
        mem[14'd2078] <= 32'h3c8dd4ab;
        mem[14'd2079] <= 32'h3c4a0677;
        mem[14'd2080] <= 32'h3c71a7a3;
        mem[14'd2081] <= 32'hbca05b3c;
        mem[14'd2082] <= 32'hbd854a4d;
        mem[14'd2083] <= 32'hbdd8def2;
        mem[14'd2084] <= 32'hbdbbf069;
        mem[14'd2085] <= 32'hbe7c0d02;
        mem[14'd2086] <= 32'hbf13d3b8;
        mem[14'd2087] <= 32'hbf05a9e6;
        mem[14'd2088] <= 32'hbca9ecd0;
        mem[14'd2089] <= 32'h3eae2cc4;
        mem[14'd2090] <= 32'h3f0ee2bc;
        mem[14'd2091] <= 32'h3ec1f45a;
        mem[14'd2092] <= 32'h3e0fc661;
        mem[14'd2093] <= 32'hbe300603;
        mem[14'd2094] <= 32'hbed2e71d;
        mem[14'd2095] <= 32'hbead5814;
        mem[14'd2096] <= 32'hbe58aa56;
        mem[14'd2097] <= 32'hbe1e7528;
        mem[14'd2098] <= 32'hbdb65879;
        mem[14'd2099] <= 32'hbd99dbbe;
        mem[14'd2100] <= 32'hbc80aeab;
        mem[14'd2101] <= 32'hbd12008e;
        mem[14'd2102] <= 32'h3c28ed06;
        mem[14'd2103] <= 32'hbb39b28c;
        mem[14'd2104] <= 32'hbb15535d;
        mem[14'd2105] <= 32'h3bcd2778;
        mem[14'd2106] <= 32'h3b989a03;
        mem[14'd2107] <= 32'hbbde829a;
        mem[14'd2108] <= 32'h3b340700;
        mem[14'd2109] <= 32'hbd869d44;
        mem[14'd2110] <= 32'hbddf8814;
        mem[14'd2111] <= 32'hbe0655f6;
        mem[14'd2112] <= 32'hbde5d82f;
        mem[14'd2113] <= 32'hbe8fc24c;
        mem[14'd2114] <= 32'hbece2b10;
        mem[14'd2115] <= 32'hbe5add1d;
        mem[14'd2116] <= 32'h3d99bf7d;
        mem[14'd2117] <= 32'h3ed8ba5c;
        mem[14'd2118] <= 32'h3f225bfa;
        mem[14'd2119] <= 32'h3e26ad37;
        mem[14'd2120] <= 32'h3de577b9;
        mem[14'd2121] <= 32'hbedb1a44;
        mem[14'd2122] <= 32'hbeefa628;
        mem[14'd2123] <= 32'hbec70758;
        mem[14'd2124] <= 32'hbe7d289c;
        mem[14'd2125] <= 32'hbe2b10da;
        mem[14'd2126] <= 32'hbdedf87f;
        mem[14'd2127] <= 32'hbd53110c;
        mem[14'd2128] <= 32'hbd46e857;
        mem[14'd2129] <= 32'hbc93d762;
        mem[14'd2130] <= 32'hbb2323a6;
        mem[14'd2131] <= 32'h3c99c4ea;
        mem[14'd2132] <= 32'hbb8fffe2;
        mem[14'd2133] <= 32'hbce1f315;
        mem[14'd2134] <= 32'hb9dc9837;
        mem[14'd2135] <= 32'hbb205c2a;
        mem[14'd2136] <= 32'hbc6d2287;
        mem[14'd2137] <= 32'hbdd6215c;
        mem[14'd2138] <= 32'hbe4cf5f6;
        mem[14'd2139] <= 32'hbe78bd5e;
        mem[14'd2140] <= 32'hbe67ef61;
        mem[14'd2141] <= 32'hbe3423f4;
        mem[14'd2142] <= 32'hbdf346fd;
        mem[14'd2143] <= 32'hbe082489;
        mem[14'd2144] <= 32'hbdc69a67;
        mem[14'd2145] <= 32'h3ec9cba0;
        mem[14'd2146] <= 32'h3f1bb75e;
        mem[14'd2147] <= 32'hbc7e0733;
        mem[14'd2148] <= 32'hbe25e1b9;
        mem[14'd2149] <= 32'hbf16fe0d;
        mem[14'd2150] <= 32'hbeea0ce5;
        mem[14'd2151] <= 32'hbeb44393;
        mem[14'd2152] <= 32'hbe7a85b5;
        mem[14'd2153] <= 32'hbe2a5360;
        mem[14'd2154] <= 32'hbdf8480f;
        mem[14'd2155] <= 32'hbde120b7;
        mem[14'd2156] <= 32'hbd695648;
        mem[14'd2157] <= 32'hbd1753c9;
        mem[14'd2158] <= 32'hbcb5905b;
        mem[14'd2159] <= 32'h3c700873;
        mem[14'd2160] <= 32'h3c7055a6;
        mem[14'd2161] <= 32'h3c151234;
        mem[14'd2162] <= 32'hbb7fcbf9;
        mem[14'd2163] <= 32'hbb806197;
        mem[14'd2164] <= 32'hbd080797;
        mem[14'd2165] <= 32'hbe2dcf36;
        mem[14'd2166] <= 32'hbeab8f0a;
        mem[14'd2167] <= 32'hbea35fbc;
        mem[14'd2168] <= 32'hbe77e5b0;
        mem[14'd2169] <= 32'hbdcd68fe;
        mem[14'd2170] <= 32'h3baff0a9;
        mem[14'd2171] <= 32'hbe279a3e;
        mem[14'd2172] <= 32'h3d68da08;
        mem[14'd2173] <= 32'h3ec9e264;
        mem[14'd2174] <= 32'h3ee52a17;
        mem[14'd2175] <= 32'hbcafa8c1;
        mem[14'd2176] <= 32'hbec0ba1d;
        mem[14'd2177] <= 32'hbf05eee1;
        mem[14'd2178] <= 32'hbeb29096;
        mem[14'd2179] <= 32'hbe6251aa;
        mem[14'd2180] <= 32'hbe2bc60e;
        mem[14'd2181] <= 32'hbe038980;
        mem[14'd2182] <= 32'hbd9de1a3;
        mem[14'd2183] <= 32'hbd82fd06;
        mem[14'd2184] <= 32'hbd3ebb4b;
        mem[14'd2185] <= 32'hbd221a72;
        mem[14'd2186] <= 32'hbc93698d;
        mem[14'd2187] <= 32'hbc342234;
        mem[14'd2188] <= 32'h3c0a8d27;
        mem[14'd2189] <= 32'hbb3710ec;
        mem[14'd2190] <= 32'hbc82c7aa;
        mem[14'd2191] <= 32'hbc50720c;
        mem[14'd2192] <= 32'hbd3bc925;
        mem[14'd2193] <= 32'hbe5ad4d8;
        mem[14'd2194] <= 32'hbeda9a30;
        mem[14'd2195] <= 32'hbeb4f9cd;
        mem[14'd2196] <= 32'hbe0b8553;
        mem[14'd2197] <= 32'hbcc01d7b;
        mem[14'd2198] <= 32'hbdfb47b0;
        mem[14'd2199] <= 32'hbe0442be;
        mem[14'd2200] <= 32'h3cec4386;
        mem[14'd2201] <= 32'h3e417612;
        mem[14'd2202] <= 32'h3e4775d0;
        mem[14'd2203] <= 32'hbe3e0ec7;
        mem[14'd2204] <= 32'hbeb27452;
        mem[14'd2205] <= 32'hbe6cdda8;
        mem[14'd2206] <= 32'hbdc3d436;
        mem[14'd2207] <= 32'hbd8bd1ab;
        mem[14'd2208] <= 32'hbcacf78d;
        mem[14'd2209] <= 32'hbd28d907;
        mem[14'd2210] <= 32'hbdbd8d7f;
        mem[14'd2211] <= 32'hbd872d1e;
        mem[14'd2212] <= 32'hbcc1b659;
        mem[14'd2213] <= 32'h3b051063;
        mem[14'd2214] <= 32'h3c3d03d0;
        mem[14'd2215] <= 32'h3bcabf23;
        mem[14'd2216] <= 32'h3c55b3ab;
        mem[14'd2217] <= 32'h3c3293da;
        mem[14'd2218] <= 32'h39b67e55;
        mem[14'd2219] <= 32'hbcb981a2;
        mem[14'd2220] <= 32'hbda6baea;
        mem[14'd2221] <= 32'hbe91cd56;
        mem[14'd2222] <= 32'hbe93440f;
        mem[14'd2223] <= 32'hbe0ab79c;
        mem[14'd2224] <= 32'hbdc517d8;
        mem[14'd2225] <= 32'hbb9e8ffd;
        mem[14'd2226] <= 32'hbd9ce7d6;
        mem[14'd2227] <= 32'hbd851a99;
        mem[14'd2228] <= 32'hbd8c98dc;
        mem[14'd2229] <= 32'h3e23931d;
        mem[14'd2230] <= 32'hbb8ddbed;
        mem[14'd2231] <= 32'hbccb2f0b;
        mem[14'd2232] <= 32'h3da77b40;
        mem[14'd2233] <= 32'hbac0de31;
        mem[14'd2234] <= 32'h3df22358;
        mem[14'd2235] <= 32'h3e00e79c;
        mem[14'd2236] <= 32'h3d923bad;
        mem[14'd2237] <= 32'hbc13ef2f;
        mem[14'd2238] <= 32'hbd81069f;
        mem[14'd2239] <= 32'hbcb0135f;
        mem[14'd2240] <= 32'h3c9d4b02;
        mem[14'd2241] <= 32'h3ce06a97;
        mem[14'd2242] <= 32'h3c7fe611;
        mem[14'd2243] <= 32'h3c3d7fd6;
        mem[14'd2244] <= 32'h3ba77da2;
        mem[14'd2245] <= 32'hbc1d2b2f;
        mem[14'd2246] <= 32'hbcbe91c0;
        mem[14'd2247] <= 32'hbcb6baec;
        mem[14'd2248] <= 32'hbd7c1ce5;
        mem[14'd2249] <= 32'hbe4169c5;
        mem[14'd2250] <= 32'hbd711811;
        mem[14'd2251] <= 32'hbbf3a27b;
        mem[14'd2252] <= 32'h3d8ce4d8;
        mem[14'd2253] <= 32'h3db57d50;
        mem[14'd2254] <= 32'h3df95992;
        mem[14'd2255] <= 32'h3e04f49b;
        mem[14'd2256] <= 32'h3d862ebf;
        mem[14'd2257] <= 32'hbcfaf99b;
        mem[14'd2258] <= 32'h3c8f4e1a;
        mem[14'd2259] <= 32'hbc87b15e;
        mem[14'd2260] <= 32'h3e3d732d;
        mem[14'd2261] <= 32'h3e738664;
        mem[14'd2262] <= 32'h3ea3925e;
        mem[14'd2263] <= 32'h3e669041;
        mem[14'd2264] <= 32'h3df47f4d;
        mem[14'd2265] <= 32'h3d5a1e8a;
        mem[14'd2266] <= 32'hbd3358c8;
        mem[14'd2267] <= 32'hbc9a66ef;
        mem[14'd2268] <= 32'hbbdd6268;
        mem[14'd2269] <= 32'h3adcd2fd;
        mem[14'd2270] <= 32'hbbcafb4d;
        mem[14'd2271] <= 32'h3b84f528;
        mem[14'd2272] <= 32'hbc4a0d80;
        mem[14'd2273] <= 32'hbb8db287;
        mem[14'd2274] <= 32'hbcca7db6;
        mem[14'd2275] <= 32'h3c2967bc;
        mem[14'd2276] <= 32'h3d289487;
        mem[14'd2277] <= 32'h3e5747a8;
        mem[14'd2278] <= 32'h3e63bdd5;
        mem[14'd2279] <= 32'h3e466eff;
        mem[14'd2280] <= 32'h3e06b8c8;
        mem[14'd2281] <= 32'h3d4c0472;
        mem[14'd2282] <= 32'h3e2de4ae;
        mem[14'd2283] <= 32'hbdb8407f;
        mem[14'd2284] <= 32'hbe1f2aac;
        mem[14'd2285] <= 32'hbe24c2b4;
        mem[14'd2286] <= 32'h3cf8b068;
        mem[14'd2287] <= 32'h3d9b84dc;
        mem[14'd2288] <= 32'h3d224f15;
        mem[14'd2289] <= 32'h3e0fd593;
        mem[14'd2290] <= 32'h3e86fc0f;
        mem[14'd2291] <= 32'h3e1e1f8e;
        mem[14'd2292] <= 32'h3e1777d3;
        mem[14'd2293] <= 32'h3da01557;
        mem[14'd2294] <= 32'hbda8bb2b;
        mem[14'd2295] <= 32'hbd8ed183;
        mem[14'd2296] <= 32'h3cdc0f7a;
        mem[14'd2297] <= 32'h3c3e1300;
        mem[14'd2298] <= 32'h3b8f6405;
        mem[14'd2299] <= 32'h3c2cbe3b;
        mem[14'd2300] <= 32'h3ca7cf55;
        mem[14'd2301] <= 32'hbbbe7ab7;
        mem[14'd2302] <= 32'h3bea95fd;
        mem[14'd2303] <= 32'hbc40128d;
        mem[14'd2304] <= 32'h3dba9a09;
        mem[14'd2305] <= 32'h3ecc9af3;
        mem[14'd2306] <= 32'h3eb035f9;
        mem[14'd2307] <= 32'h3e2a7f08;
        mem[14'd2308] <= 32'h3da03d89;
        mem[14'd2309] <= 32'h3d8100b1;
        mem[14'd2310] <= 32'hbdd729a2;
        mem[14'd2311] <= 32'hbe995cfd;
        mem[14'd2312] <= 32'hbedceded;
        mem[14'd2313] <= 32'hbeac2bfe;
        mem[14'd2314] <= 32'hbdb1b185;
        mem[14'd2315] <= 32'hbc81ff45;
        mem[14'd2316] <= 32'h3d081aa0;
        mem[14'd2317] <= 32'h3e80834c;
        mem[14'd2318] <= 32'h3e7e4624;
        mem[14'd2319] <= 32'h3e26b127;
        mem[14'd2320] <= 32'h3de1ef9e;
        mem[14'd2321] <= 32'hbca9ea07;
        mem[14'd2322] <= 32'hbe01bb88;
        mem[14'd2323] <= 32'hbd801640;
        mem[14'd2324] <= 32'hbb7d0b2b;
        mem[14'd2325] <= 32'h3c61b4aa;
        mem[14'd2326] <= 32'h39e08f10;
        mem[14'd2327] <= 32'hbabaabb8;
        mem[14'd2328] <= 32'hbc237567;
        mem[14'd2329] <= 32'hbb81afbc;
        mem[14'd2330] <= 32'hbaf0025d;
        mem[14'd2331] <= 32'hbc79a15d;
        mem[14'd2332] <= 32'h3cf1e1c5;
        mem[14'd2333] <= 32'h3e6c88b9;
        mem[14'd2334] <= 32'h3e7cce40;
        mem[14'd2335] <= 32'h3dc15329;
        mem[14'd2336] <= 32'hbcf88b83;
        mem[14'd2337] <= 32'hbd1709b1;
        mem[14'd2338] <= 32'hbdc82b3f;
        mem[14'd2339] <= 32'hbe1839ce;
        mem[14'd2340] <= 32'hbcb65660;
        mem[14'd2341] <= 32'hbe08aa58;
        mem[14'd2342] <= 32'hbe2ede14;
        mem[14'd2343] <= 32'h3c4cc889;
        mem[14'd2344] <= 32'h3dac8ccb;
        mem[14'd2345] <= 32'h3e4d3609;
        mem[14'd2346] <= 32'h3d85b66e;
        mem[14'd2347] <= 32'h3d5d627f;
        mem[14'd2348] <= 32'hbc4e133a;
        mem[14'd2349] <= 32'hbdaf105e;
        mem[14'd2350] <= 32'hbd96b6b1;
        mem[14'd2351] <= 32'hbd3d7c5a;
        mem[14'd2352] <= 32'h3a3cf3ef;
        mem[14'd2353] <= 32'h3c13e888;
        mem[14'd2354] <= 32'h3c19a207;
        mem[14'd2355] <= 32'hbc603041;
        mem[14'd2356] <= 32'h3b13c004;
        mem[14'd2357] <= 32'hbbc737fc;
        mem[14'd2358] <= 32'h3ae7267d;
        mem[14'd2359] <= 32'hbccaa91e;
        mem[14'd2360] <= 32'hbcfcc7f2;
        mem[14'd2361] <= 32'h3c8db97e;
        mem[14'd2362] <= 32'h3cfe08e0;
        mem[14'd2363] <= 32'hbd9c562e;
        mem[14'd2364] <= 32'hbe44ce41;
        mem[14'd2365] <= 32'hbe2e44be;
        mem[14'd2366] <= 32'hbe666b8c;
        mem[14'd2367] <= 32'hbe91366e;
        mem[14'd2368] <= 32'hbe7b416b;
        mem[14'd2369] <= 32'hbe982085;
        mem[14'd2370] <= 32'hbe983054;
        mem[14'd2371] <= 32'hbe7be079;
        mem[14'd2372] <= 32'hbe992bfa;
        mem[14'd2373] <= 32'hbdac271f;
        mem[14'd2374] <= 32'hbba9f926;
        mem[14'd2375] <= 32'h3ca51444;
        mem[14'd2376] <= 32'hbcc10c16;
        mem[14'd2377] <= 32'hbcd7280f;
        mem[14'd2378] <= 32'hbd2127e4;
        mem[14'd2379] <= 32'hbc371ddb;
        mem[14'd2380] <= 32'hbbf470ac;
        mem[14'd2381] <= 32'h3a9aa95f;
        mem[14'd2382] <= 32'hbbcc00de;
        mem[14'd2383] <= 32'h3c366507;
        mem[14'd2384] <= 32'hbbc6c8ca;
        mem[14'd2385] <= 32'h3c8fa5c3;
        mem[14'd2386] <= 32'h3c11984e;
        mem[14'd2387] <= 32'hbb449e01;
        mem[14'd2388] <= 32'hbd0f0cfd;
        mem[14'd2389] <= 32'hbd568732;
        mem[14'd2390] <= 32'hbd8e2839;
        mem[14'd2391] <= 32'hbdc69f3b;
        mem[14'd2392] <= 32'hbdcf3866;
        mem[14'd2393] <= 32'hbe232969;
        mem[14'd2394] <= 32'hbe9ea659;
        mem[14'd2395] <= 32'hbe919606;
        mem[14'd2396] <= 32'hbe50d297;
        mem[14'd2397] <= 32'hbe82c7af;
        mem[14'd2398] <= 32'hbe82c559;
        mem[14'd2399] <= 32'hbe86d258;
        mem[14'd2400] <= 32'hbe5866d0;
        mem[14'd2401] <= 32'hbe0a1647;
        mem[14'd2402] <= 32'hbd35f875;
        mem[14'd2403] <= 32'hbd332565;
        mem[14'd2404] <= 32'hbc4b2a0c;
        mem[14'd2405] <= 32'h3b29576d;
        mem[14'd2406] <= 32'h3b6e3cef;
        mem[14'd2407] <= 32'hbac5237b;
        mem[14'd2408] <= 32'h3bbdfb17;
        mem[14'd2409] <= 32'h3aa7ec94;
        mem[14'd2410] <= 32'h3bd68af8;
        mem[14'd2411] <= 32'h3c58d4ce;
        mem[14'd2412] <= 32'h3bbad315;
        mem[14'd2413] <= 32'h3af876b5;
        mem[14'd2414] <= 32'h3c5d1712;
        mem[14'd2415] <= 32'h3b03bf65;
        mem[14'd2416] <= 32'hbbe992a6;
        mem[14'd2417] <= 32'hbb9f6568;
        mem[14'd2418] <= 32'hbc50af6e;
        mem[14'd2419] <= 32'hbc7c07cb;
        mem[14'd2420] <= 32'hbca08ffb;
        mem[14'd2421] <= 32'hbc849c98;
        mem[14'd2422] <= 32'hbd5ce089;
        mem[14'd2423] <= 32'hbd3a3c93;
        mem[14'd2424] <= 32'hbd81f70b;
        mem[14'd2425] <= 32'hbd7f3146;
        mem[14'd2426] <= 32'hbd81481a;
        mem[14'd2427] <= 32'hbd5ce986;
        mem[14'd2428] <= 32'hbd4662da;
        mem[14'd2429] <= 32'hbc80a213;
        mem[14'd2430] <= 32'hbd26e2fe;
        mem[14'd2431] <= 32'h3a845980;
        mem[14'd2432] <= 32'h3b7d3a4a;
        mem[14'd2433] <= 32'hbc169991;
        mem[14'd2434] <= 32'hbbbae6f8;
        mem[14'd2435] <= 32'h3ba1b623;
        mem[14'd2436] <= 32'h3c5308ec;
        mem[14'd2437] <= 32'hba862224;
        mem[14'd2438] <= 32'hbb8b0566;
        mem[14'd2439] <= 32'hbbeb6802;
        mem[14'd2440] <= 32'h3c97f50d;
        mem[14'd2441] <= 32'h3c1c13b3;
        mem[14'd2442] <= 32'h3c1718cd;
        mem[14'd2443] <= 32'hbc1867e3;
        mem[14'd2444] <= 32'h3a954148;
        mem[14'd2445] <= 32'hbc5ffe37;
        mem[14'd2446] <= 32'h3bb63bc8;
        mem[14'd2447] <= 32'hbc4aa47e;
        mem[14'd2448] <= 32'hbb3a0105;
        mem[14'd2449] <= 32'h3b907dcd;
        mem[14'd2450] <= 32'h3c5a95a8;
        mem[14'd2451] <= 32'hba9f5851;
        mem[14'd2452] <= 32'hbc3688d5;
        mem[14'd2453] <= 32'h3bd1b031;
        mem[14'd2454] <= 32'h3c65e402;
        mem[14'd2455] <= 32'h3b8e0c3a;
        mem[14'd2456] <= 32'h3c89ccae;
        mem[14'd2457] <= 32'h3bf6a040;
        mem[14'd2458] <= 32'hba9e5286;
        mem[14'd2459] <= 32'hba1556ef;
        mem[14'd2460] <= 32'hbc8755a4;
        mem[14'd2461] <= 32'hbb7f3d37;
        mem[14'd2462] <= 32'h3bca9e10;
        mem[14'd2463] <= 32'hbb280114;
        mem[14'd2464] <= 32'hbbc92e8d;
        mem[14'd2465] <= 32'hbca81907;
        mem[14'd2466] <= 32'hbc2b429b;
        mem[14'd2467] <= 32'h3bef8067;
        mem[14'd2468] <= 32'h3bc00a82;
        mem[14'd2469] <= 32'hbc936f4f;
        mem[14'd2470] <= 32'h3a2ad45b;
        mem[14'd2471] <= 32'hbc15da8b;
        mem[14'd2472] <= 32'h3c9ec607;
        mem[14'd2473] <= 32'hbc8d5661;
        mem[14'd2474] <= 32'h394ba28b;
        mem[14'd2475] <= 32'hbbb2f40e;
        mem[14'd2476] <= 32'hbc875e75;
        mem[14'd2477] <= 32'h3c3022ca;
        mem[14'd2478] <= 32'h3b5e1f7d;
        mem[14'd2479] <= 32'hbbc23577;
        mem[14'd2480] <= 32'hbb84a121;
        mem[14'd2481] <= 32'h3c30e39a;
        mem[14'd2482] <= 32'h3b257e19;
        mem[14'd2483] <= 32'h3c03d81a;
        mem[14'd2484] <= 32'hbc97eb8f;
        mem[14'd2485] <= 32'h3be00ee7;
        mem[14'd2486] <= 32'hbb3cb76f;
        mem[14'd2487] <= 32'hbc8140e4;
        mem[14'd2488] <= 32'hbc4ec784;
        mem[14'd2489] <= 32'hbbfc06b8;
        mem[14'd2490] <= 32'h3bbb1d69;
        mem[14'd2491] <= 32'hbb8f641b;
        mem[14'd2492] <= 32'hb8b73112;
        mem[14'd2493] <= 32'hbb980b7d;
        mem[14'd2494] <= 32'hbc365820;
        mem[14'd2495] <= 32'h3c01dab9;
        mem[14'd2496] <= 32'hbbf3eaf3;
        mem[14'd2497] <= 32'h3c51d480;
        mem[14'd2498] <= 32'h3c6a877d;
        mem[14'd2499] <= 32'hbc237be4;
        mem[14'd2500] <= 32'h3c16ef1f;
        mem[14'd2501] <= 32'h3cbfca75;
        mem[14'd2502] <= 32'h3be40fba;
        mem[14'd2503] <= 32'hbbddee14;
        mem[14'd2504] <= 32'hbbede789;
        mem[14'd2505] <= 32'hbb6a7ec1;
        mem[14'd2506] <= 32'hbcbb828c;
        mem[14'd2507] <= 32'hbbd86c38;
        mem[14'd2508] <= 32'hba09a102;
        mem[14'd2509] <= 32'hbc8b131d;
        mem[14'd2510] <= 32'hbc0ce973;
        mem[14'd2511] <= 32'h3c98391c;
        mem[14'd2512] <= 32'h3d44d90b;
        mem[14'd2513] <= 32'h3bd752cd;
        mem[14'd2514] <= 32'h3a94968a;
        mem[14'd2515] <= 32'hbbddf336;
        mem[14'd2516] <= 32'h3ba35a84;
        mem[14'd2517] <= 32'h3b32e7ad;
        mem[14'd2518] <= 32'h3ab2a177;
        mem[14'd2519] <= 32'hbc165cc3;
        mem[14'd2520] <= 32'h3b1a48c6;
        mem[14'd2521] <= 32'hba872a60;
        mem[14'd2522] <= 32'hba6ea733;
        mem[14'd2523] <= 32'hbaecc981;
        mem[14'd2524] <= 32'h3bf0539e;
        mem[14'd2525] <= 32'hbc08257d;
        mem[14'd2526] <= 32'h3bcd883e;
        mem[14'd2527] <= 32'h3b457dfe;
        mem[14'd2528] <= 32'hbb99c947;
        mem[14'd2529] <= 32'hbc111b60;
        mem[14'd2530] <= 32'hbc301da3;
        mem[14'd2531] <= 32'h3b53bec0;
        mem[14'd2532] <= 32'hbb24a99d;
        mem[14'd2533] <= 32'h3c4e3111;
        mem[14'd2534] <= 32'h3d01ddca;
        mem[14'd2535] <= 32'h3d0fc90f;
        mem[14'd2536] <= 32'h3d6bd7fd;
        mem[14'd2537] <= 32'h3d47a4f6;
        mem[14'd2538] <= 32'h3d39a7df;
        mem[14'd2539] <= 32'h3d959ee5;
        mem[14'd2540] <= 32'h3da9b488;
        mem[14'd2541] <= 32'h3d091757;
        mem[14'd2542] <= 32'hbd0b3951;
        mem[14'd2543] <= 32'hbd5cbcde;
        mem[14'd2544] <= 32'hbd1fc9df;
        mem[14'd2545] <= 32'hbd1f44ea;
        mem[14'd2546] <= 32'hbcda264f;
        mem[14'd2547] <= 32'hbc96a9d1;
        mem[14'd2548] <= 32'h3cfb9ef6;
        mem[14'd2549] <= 32'h3c83adfc;
        mem[14'd2550] <= 32'hbbf608fe;
        mem[14'd2551] <= 32'hbc7108a5;
        mem[14'd2552] <= 32'hbc87f7d1;
        mem[14'd2553] <= 32'h3c8ce98d;
        mem[14'd2554] <= 32'h3bcc3256;
        mem[14'd2555] <= 32'hb9f54fc0;
        mem[14'd2556] <= 32'hbbc7ff54;
        mem[14'd2557] <= 32'h3acf4dbb;
        mem[14'd2558] <= 32'h3ac1a64a;
        mem[14'd2559] <= 32'h3c5043fb;
        mem[14'd2560] <= 32'h3d922027;
        mem[14'd2561] <= 32'h3e552bb5;
        mem[14'd2562] <= 32'h3e83a3af;
        mem[14'd2563] <= 32'h3e96d007;
        mem[14'd2564] <= 32'h3ea5451c;
        mem[14'd2565] <= 32'h3eb1ccb6;
        mem[14'd2566] <= 32'h3e799df5;
        mem[14'd2567] <= 32'h3e1cb13d;
        mem[14'd2568] <= 32'h3e4134f9;
        mem[14'd2569] <= 32'h3db3c178;
        mem[14'd2570] <= 32'hbd9e2beb;
        mem[14'd2571] <= 32'hbdfd5ada;
        mem[14'd2572] <= 32'hbe0f86b1;
        mem[14'd2573] <= 32'hbdcc7bfe;
        mem[14'd2574] <= 32'hbdd20ca8;
        mem[14'd2575] <= 32'hbd5f769a;
        mem[14'd2576] <= 32'hbc9ed27f;
        mem[14'd2577] <= 32'h3c02197b;
        mem[14'd2578] <= 32'h3b38066c;
        mem[14'd2579] <= 32'h3c233cb9;
        mem[14'd2580] <= 32'hbbe93410;
        mem[14'd2581] <= 32'h3c6eac72;
        mem[14'd2582] <= 32'h3ba11d9b;
        mem[14'd2583] <= 32'hbc0ff50c;
        mem[14'd2584] <= 32'hbccd5ab1;
        mem[14'd2585] <= 32'h3c1afd5d;
        mem[14'd2586] <= 32'h3d8040b9;
        mem[14'd2587] <= 32'h3d942543;
        mem[14'd2588] <= 32'h3de829f1;
        mem[14'd2589] <= 32'h3e8d92f3;
        mem[14'd2590] <= 32'h3e819243;
        mem[14'd2591] <= 32'h3e93e435;
        mem[14'd2592] <= 32'h3e8fcca9;
        mem[14'd2593] <= 32'h3e475700;
        mem[14'd2594] <= 32'h3e6848fb;
        mem[14'd2595] <= 32'h3ddfb536;
        mem[14'd2596] <= 32'h3dad185a;
        mem[14'd2597] <= 32'h3db0717c;
        mem[14'd2598] <= 32'hbcc43094;
        mem[14'd2599] <= 32'hbde527ee;
        mem[14'd2600] <= 32'hbe0364e7;
        mem[14'd2601] <= 32'hbe731851;
        mem[14'd2602] <= 32'hbe83e425;
        mem[14'd2603] <= 32'hbe395fcc;
        mem[14'd2604] <= 32'hbdaf0a67;
        mem[14'd2605] <= 32'hbc93fadc;
        mem[14'd2606] <= 32'hbbae2640;
        mem[14'd2607] <= 32'h3b4e3a29;
        mem[14'd2608] <= 32'hbb91a140;
        mem[14'd2609] <= 32'hbc3d93c5;
        mem[14'd2610] <= 32'hbbc0f630;
        mem[14'd2611] <= 32'hbc8acbb5;
        mem[14'd2612] <= 32'hb9317fec;
        mem[14'd2613] <= 32'h3d57a9ba;
        mem[14'd2614] <= 32'h3d90b1c8;
        mem[14'd2615] <= 32'h3decb854;
        mem[14'd2616] <= 32'h3e4f7bcc;
        mem[14'd2617] <= 32'h3e42b1a2;
        mem[14'd2618] <= 32'h3e42000e;
        mem[14'd2619] <= 32'h3e84ca94;
        mem[14'd2620] <= 32'h3e5aa7b1;
        mem[14'd2621] <= 32'h3e566068;
        mem[14'd2622] <= 32'h3e285375;
        mem[14'd2623] <= 32'h3e302ab2;
        mem[14'd2624] <= 32'h3e9007c4;
        mem[14'd2625] <= 32'h3e5caa40;
        mem[14'd2626] <= 32'h3e0b016f;
        mem[14'd2627] <= 32'h3ccb9a58;
        mem[14'd2628] <= 32'hbc99a544;
        mem[14'd2629] <= 32'hbd2e9872;
        mem[14'd2630] <= 32'hbe17689d;
        mem[14'd2631] <= 32'hbe5039e7;
        mem[14'd2632] <= 32'hbe1735e1;
        mem[14'd2633] <= 32'hbd0bf3e0;
        mem[14'd2634] <= 32'hbc951fc4;
        mem[14'd2635] <= 32'h3c0a5a42;
        mem[14'd2636] <= 32'h3b38f65e;
        mem[14'd2637] <= 32'hbc63d33d;
        mem[14'd2638] <= 32'hbcf60990;
        mem[14'd2639] <= 32'h3c812d5d;
        mem[14'd2640] <= 32'h3d9a9293;
        mem[14'd2641] <= 32'h3dc81343;
        mem[14'd2642] <= 32'h3e1165c6;
        mem[14'd2643] <= 32'h3e2e1f7d;
        mem[14'd2644] <= 32'h3e02edae;
        mem[14'd2645] <= 32'h3e1b1602;
        mem[14'd2646] <= 32'h3e10e38a;
        mem[14'd2647] <= 32'h3d064cd5;
        mem[14'd2648] <= 32'h3cae60bf;
        mem[14'd2649] <= 32'h3db43592;
        mem[14'd2650] <= 32'h3d99193a;
        mem[14'd2651] <= 32'h3dcaff1a;
        mem[14'd2652] <= 32'h3deca6a4;
        mem[14'd2653] <= 32'h3d121a33;
        mem[14'd2654] <= 32'h3ccc4f48;
        mem[14'd2655] <= 32'hbd8d98f3;
        mem[14'd2656] <= 32'hbda80579;
        mem[14'd2657] <= 32'hbda29432;
        mem[14'd2658] <= 32'hbe3d469b;
        mem[14'd2659] <= 32'hbea9063f;
        mem[14'd2660] <= 32'hbe308a82;
        mem[14'd2661] <= 32'hbd64e9d4;
        mem[14'd2662] <= 32'hbcabf46f;
        mem[14'd2663] <= 32'hbc89877c;
        mem[14'd2664] <= 32'h3c16b0db;
        mem[14'd2665] <= 32'h3c16b24d;
        mem[14'd2666] <= 32'hbb557685;
        mem[14'd2667] <= 32'h3cefdfe5;
        mem[14'd2668] <= 32'h3e186958;
        mem[14'd2669] <= 32'h3e20feac;
        mem[14'd2670] <= 32'h3e5ffaeb;
        mem[14'd2671] <= 32'h3db20fa3;
        mem[14'd2672] <= 32'h3e0962d7;
        mem[14'd2673] <= 32'h3cef5427;
        mem[14'd2674] <= 32'hbc7d2fee;
        mem[14'd2675] <= 32'h3dc5486c;
        mem[14'd2676] <= 32'hbc65a4e4;
        mem[14'd2677] <= 32'h3e1b591c;
        mem[14'd2678] <= 32'h3d210b1d;
        mem[14'd2679] <= 32'hbd9560a3;
        mem[14'd2680] <= 32'hbc89388b;
        mem[14'd2681] <= 32'hbe711538;
        mem[14'd2682] <= 32'hbdaa30e3;
        mem[14'd2683] <= 32'hbd8cdb5f;
        mem[14'd2684] <= 32'hbdea5182;
        mem[14'd2685] <= 32'h3b8834fa;
        mem[14'd2686] <= 32'h3c4149cb;
        mem[14'd2687] <= 32'hbeae2e7a;
        mem[14'd2688] <= 32'hbe6c7836;
        mem[14'd2689] <= 32'hbda21aca;
        mem[14'd2690] <= 32'hbc826a72;
        mem[14'd2691] <= 32'h3b074b93;
        mem[14'd2692] <= 32'hbbc7687f;
        mem[14'd2693] <= 32'hbc02225e;
        mem[14'd2694] <= 32'h3c377d53;
        mem[14'd2695] <= 32'h3d066153;
        mem[14'd2696] <= 32'h3e38968a;
        mem[14'd2697] <= 32'h3e1a7130;
        mem[14'd2698] <= 32'h3dc75b4d;
        mem[14'd2699] <= 32'h3da1ef13;
        mem[14'd2700] <= 32'h3d741387;
        mem[14'd2701] <= 32'h3cdfff85;
        mem[14'd2702] <= 32'h3e5fced0;
        mem[14'd2703] <= 32'h3dfc85d0;
        mem[14'd2704] <= 32'hbc9d4c7e;
        mem[14'd2705] <= 32'hbcbaaedf;
        mem[14'd2706] <= 32'h3d85a97c;
        mem[14'd2707] <= 32'h3d08e3b4;
        mem[14'd2708] <= 32'hbd53d3d4;
        mem[14'd2709] <= 32'hbc94294b;
        mem[14'd2710] <= 32'hbe08e476;
        mem[14'd2711] <= 32'h3dc4a009;
        mem[14'd2712] <= 32'h3d068cbd;
        mem[14'd2713] <= 32'hbccd861d;
        mem[14'd2714] <= 32'hbcbe082e;
        mem[14'd2715] <= 32'hbe12d557;
        mem[14'd2716] <= 32'hbe8998fd;
        mem[14'd2717] <= 32'hbdd1241b;
        mem[14'd2718] <= 32'hbbcc84af;
        mem[14'd2719] <= 32'hbc923bba;
        mem[14'd2720] <= 32'hbb4fdfa5;
        mem[14'd2721] <= 32'hbc8c0852;
        mem[14'd2722] <= 32'hbc5bdc5e;
        mem[14'd2723] <= 32'h3cf0ccfa;
        mem[14'd2724] <= 32'h3e010e23;
        mem[14'd2725] <= 32'h3e55426c;
        mem[14'd2726] <= 32'h3d60ccf0;
        mem[14'd2727] <= 32'h3bb28f82;
        mem[14'd2728] <= 32'hbd2cfd08;
        mem[14'd2729] <= 32'h3df3a620;
        mem[14'd2730] <= 32'h3e39343b;
        mem[14'd2731] <= 32'h3d40083d;
        mem[14'd2732] <= 32'h3d13a2c0;
        mem[14'd2733] <= 32'h3db038a5;
        mem[14'd2734] <= 32'h3e109100;
        mem[14'd2735] <= 32'h3e37fff3;
        mem[14'd2736] <= 32'h3dfd64d9;
        mem[14'd2737] <= 32'h3cdf9053;
        mem[14'd2738] <= 32'h3da46f3e;
        mem[14'd2739] <= 32'h3cbada61;
        mem[14'd2740] <= 32'hbbf82745;
        mem[14'd2741] <= 32'hbdb4e106;
        mem[14'd2742] <= 32'hbb71b25c;
        mem[14'd2743] <= 32'hbdfd8170;
        mem[14'd2744] <= 32'hbe74ca5b;
        mem[14'd2745] <= 32'hbdb77772;
        mem[14'd2746] <= 32'hbcd94d33;
        mem[14'd2747] <= 32'h3b86a59d;
        mem[14'd2748] <= 32'hbc50295c;
        mem[14'd2749] <= 32'h3c21e0b2;
        mem[14'd2750] <= 32'hbbec74a1;
        mem[14'd2751] <= 32'h3d2f008b;
        mem[14'd2752] <= 32'h3ca0e312;
        mem[14'd2753] <= 32'h3df91f62;
        mem[14'd2754] <= 32'h3e1589dd;
        mem[14'd2755] <= 32'hbd838219;
        mem[14'd2756] <= 32'hbd2e5242;
        mem[14'd2757] <= 32'hbdfaef9e;
        mem[14'd2758] <= 32'hbdcbdfff;
        mem[14'd2759] <= 32'hbd924e34;
        mem[14'd2760] <= 32'hbdf8a3ec;
        mem[14'd2761] <= 32'hbe799166;
        mem[14'd2762] <= 32'hbd8658a8;
        mem[14'd2763] <= 32'hbdcb8840;
        mem[14'd2764] <= 32'h3c4f1864;
        mem[14'd2765] <= 32'h3de58a55;
        mem[14'd2766] <= 32'h3d5b8acc;
        mem[14'd2767] <= 32'hbd2899c6;
        mem[14'd2768] <= 32'hbbc5d91f;
        mem[14'd2769] <= 32'hbd84879c;
        mem[14'd2770] <= 32'hbcfcb3ea;
        mem[14'd2771] <= 32'hbdfc96dc;
        mem[14'd2772] <= 32'hbe2862e0;
        mem[14'd2773] <= 32'hbd443104;
        mem[14'd2774] <= 32'h3c353211;
        mem[14'd2775] <= 32'h3c26660e;
        mem[14'd2776] <= 32'h3be7308f;
        mem[14'd2777] <= 32'hbb37f184;
        mem[14'd2778] <= 32'h3c588532;
        mem[14'd2779] <= 32'hbc91ac47;
        mem[14'd2780] <= 32'hbd895b03;
        mem[14'd2781] <= 32'hbdbdcff9;
        mem[14'd2782] <= 32'hbe4fb63f;
        mem[14'd2783] <= 32'hbeb457d5;
        mem[14'd2784] <= 32'hbec688d2;
        mem[14'd2785] <= 32'hbef4a2ba;
        mem[14'd2786] <= 32'hbf216732;
        mem[14'd2787] <= 32'hbf13b6e3;
        mem[14'd2788] <= 32'hbf22cc88;
        mem[14'd2789] <= 32'hbf3e149a;
        mem[14'd2790] <= 32'hbf05a88f;
        mem[14'd2791] <= 32'hbebe0b60;
        mem[14'd2792] <= 32'hbe159c5b;
        mem[14'd2793] <= 32'hbe819e7e;
        mem[14'd2794] <= 32'hbdd1e7f1;
        mem[14'd2795] <= 32'h3dc705b5;
        mem[14'd2796] <= 32'hbd8c2dbf;
        mem[14'd2797] <= 32'hbd34274a;
        mem[14'd2798] <= 32'hbd8c5882;
        mem[14'd2799] <= 32'hbde95dbd;
        mem[14'd2800] <= 32'hbd675c71;
        mem[14'd2801] <= 32'h3d692191;
        mem[14'd2802] <= 32'h3c5b87c6;
        mem[14'd2803] <= 32'h3c028eb5;
        mem[14'd2804] <= 32'h3cae4eca;
        mem[14'd2805] <= 32'hbb977152;
        mem[14'd2806] <= 32'hbcab0f6b;
        mem[14'd2807] <= 32'hbda28532;
        mem[14'd2808] <= 32'hbe28130e;
        mem[14'd2809] <= 32'hbecd4b2d;
        mem[14'd2810] <= 32'hbf2b7bbe;
        mem[14'd2811] <= 32'hbf4b4953;
        mem[14'd2812] <= 32'hbf03d81d;
        mem[14'd2813] <= 32'hbf02cb95;
        mem[14'd2814] <= 32'hbf0d8d9a;
        mem[14'd2815] <= 32'hbf044926;
        mem[14'd2816] <= 32'hbf051b53;
        mem[14'd2817] <= 32'hbeee5d17;
        mem[14'd2818] <= 32'hbec55a19;
        mem[14'd2819] <= 32'hbed36add;
        mem[14'd2820] <= 32'hbe8ce832;
        mem[14'd2821] <= 32'hbe9112e6;
        mem[14'd2822] <= 32'hbe365a57;
        mem[14'd2823] <= 32'h3da3abfc;
        mem[14'd2824] <= 32'hbd20aafb;
        mem[14'd2825] <= 32'hbca52ddb;
        mem[14'd2826] <= 32'hbde75837;
        mem[14'd2827] <= 32'hbe661cdb;
        mem[14'd2828] <= 32'h3ce5b126;
        mem[14'd2829] <= 32'h3e32b274;
        mem[14'd2830] <= 32'h3db000f5;
        mem[14'd2831] <= 32'h3c9292c4;
        mem[14'd2832] <= 32'hbc3c22b8;
        mem[14'd2833] <= 32'h3c0e61c0;
        mem[14'd2834] <= 32'hbbbcacd4;
        mem[14'd2835] <= 32'hbd69c003;
        mem[14'd2836] <= 32'hbe91c127;
        mem[14'd2837] <= 32'hbf194008;
        mem[14'd2838] <= 32'hbf449107;
        mem[14'd2839] <= 32'hbf23f004;
        mem[14'd2840] <= 32'hbec0f81f;
        mem[14'd2841] <= 32'hbe8dcd99;
        mem[14'd2842] <= 32'hbe2a882a;
        mem[14'd2843] <= 32'hbce09ebc;
        mem[14'd2844] <= 32'hbd9e0ab7;
        mem[14'd2845] <= 32'h3d5bc711;
        mem[14'd2846] <= 32'hbcea716d;
        mem[14'd2847] <= 32'hbe87746a;
        mem[14'd2848] <= 32'hbe578dd7;
        mem[14'd2849] <= 32'hbdf17f5b;
        mem[14'd2850] <= 32'hbe12f27b;
        mem[14'd2851] <= 32'hbddb329c;
        mem[14'd2852] <= 32'hbdb6ad09;
        mem[14'd2853] <= 32'hbc776968;
        mem[14'd2854] <= 32'hbdbad427;
        mem[14'd2855] <= 32'hbd90f3d9;
        mem[14'd2856] <= 32'h3e587b77;
        mem[14'd2857] <= 32'h3e8ebc0a;
        mem[14'd2858] <= 32'h3e41b5d7;
        mem[14'd2859] <= 32'h3d2936a4;
        mem[14'd2860] <= 32'h3ae6428b;
        mem[14'd2861] <= 32'hbb64a203;
        mem[14'd2862] <= 32'hbbb6c84b;
        mem[14'd2863] <= 32'hbd83b2ee;
        mem[14'd2864] <= 32'hbe50b52a;
        mem[14'd2865] <= 32'hbee44465;
        mem[14'd2866] <= 32'hbea475f0;
        mem[14'd2867] <= 32'hbdc0c09a;
        mem[14'd2868] <= 32'hbda98888;
        mem[14'd2869] <= 32'hbda59fcb;
        mem[14'd2870] <= 32'hbc0a0eea;
        mem[14'd2871] <= 32'h3d28a958;
        mem[14'd2872] <= 32'h3bd96d61;
        mem[14'd2873] <= 32'h3e6b236d;
        mem[14'd2874] <= 32'h3d8e5f41;
        mem[14'd2875] <= 32'hbddb4b31;
        mem[14'd2876] <= 32'hbdf080ee;
        mem[14'd2877] <= 32'hbe45480b;
        mem[14'd2878] <= 32'hbd120feb;
        mem[14'd2879] <= 32'hbdd23779;
        mem[14'd2880] <= 32'hbcd67e51;
        mem[14'd2881] <= 32'hbe05346f;
        mem[14'd2882] <= 32'hbdc9ed80;
        mem[14'd2883] <= 32'h3d3396d4;
        mem[14'd2884] <= 32'h3e79cb06;
        mem[14'd2885] <= 32'h3e9798b1;
        mem[14'd2886] <= 32'h3e460d0d;
        mem[14'd2887] <= 32'h3b16f38e;
        mem[14'd2888] <= 32'hbc3fcb6f;
        mem[14'd2889] <= 32'hbc2c5b28;
        mem[14'd2890] <= 32'hbcb5a966;
        mem[14'd2891] <= 32'h3d4ea89b;
        mem[14'd2892] <= 32'h3d594b40;
        mem[14'd2893] <= 32'h3db2d721;
        mem[14'd2894] <= 32'h3e3008f8;
        mem[14'd2895] <= 32'h3dafdc56;
        mem[14'd2896] <= 32'h3d05f7d8;
        mem[14'd2897] <= 32'h3d262467;
        mem[14'd2898] <= 32'h3cba0458;
        mem[14'd2899] <= 32'hbbeffa6c;
        mem[14'd2900] <= 32'hbce3f369;
        mem[14'd2901] <= 32'h3e537b12;
        mem[14'd2902] <= 32'h3db970c0;
        mem[14'd2903] <= 32'h3c7f74a4;
        mem[14'd2904] <= 32'hbcea9298;
        mem[14'd2905] <= 32'hbdfc499a;
        mem[14'd2906] <= 32'hbe018788;
        mem[14'd2907] <= 32'hbd51ee68;
        mem[14'd2908] <= 32'hbe415840;
        mem[14'd2909] <= 32'hbdecf725;
        mem[14'd2910] <= 32'hbe3f4232;
        mem[14'd2911] <= 32'hbc7d532c;
        mem[14'd2912] <= 32'h3eb9a266;
        mem[14'd2913] <= 32'h3ee28319;
        mem[14'd2914] <= 32'h3e53b195;
        mem[14'd2915] <= 32'h3c95b3b7;
        mem[14'd2916] <= 32'hbc4a47b8;
        mem[14'd2917] <= 32'hbc4b712c;
        mem[14'd2918] <= 32'h3ab8be6b;
        mem[14'd2919] <= 32'h3e25d748;
        mem[14'd2920] <= 32'h3e72ba31;
        mem[14'd2921] <= 32'h3e783f65;
        mem[14'd2922] <= 32'h3e8d7688;
        mem[14'd2923] <= 32'h3da2b8b4;
        mem[14'd2924] <= 32'hbdacd7cc;
        mem[14'd2925] <= 32'h3dfd457b;
        mem[14'd2926] <= 32'h3e172110;
        mem[14'd2927] <= 32'h3e280ef4;
        mem[14'd2928] <= 32'h3e995da1;
        mem[14'd2929] <= 32'h3ea8c0af;
        mem[14'd2930] <= 32'h3e118b41;
        mem[14'd2931] <= 32'hbc03027f;
        mem[14'd2932] <= 32'h3e090100;
        mem[14'd2933] <= 32'h3e39c05a;
        mem[14'd2934] <= 32'h3cc54f29;
        mem[14'd2935] <= 32'hbaa4b2fe;
        mem[14'd2936] <= 32'hbdcd7f0c;
        mem[14'd2937] <= 32'h3e3f6e77;
        mem[14'd2938] <= 32'h3df38f3e;
        mem[14'd2939] <= 32'h3e1ac06f;
        mem[14'd2940] <= 32'h3ee1ff04;
        mem[14'd2941] <= 32'h3f1db6af;
        mem[14'd2942] <= 32'h3e90081a;
        mem[14'd2943] <= 32'h3d1202f7;
        mem[14'd2944] <= 32'hbc2af1c5;
        mem[14'd2945] <= 32'hba681ea7;
        mem[14'd2946] <= 32'h3c37feb4;
        mem[14'd2947] <= 32'h3e2227dd;
        mem[14'd2948] <= 32'h3ea6de0f;
        mem[14'd2949] <= 32'h3e9ee4d4;
        mem[14'd2950] <= 32'h3e73a446;
        mem[14'd2951] <= 32'h3de12ac6;
        mem[14'd2952] <= 32'h3d91e8fe;
        mem[14'd2953] <= 32'h3e24711f;
        mem[14'd2954] <= 32'h3e8bbab7;
        mem[14'd2955] <= 32'h3e9cd7fd;
        mem[14'd2956] <= 32'h3eaa954a;
        mem[14'd2957] <= 32'h3e8a91d2;
        mem[14'd2958] <= 32'h3d48cfa8;
        mem[14'd2959] <= 32'h3dbace58;
        mem[14'd2960] <= 32'h3d082720;
        mem[14'd2961] <= 32'hbd17b35d;
        mem[14'd2962] <= 32'h3d2da7a8;
        mem[14'd2963] <= 32'h3c7ee0a4;
        mem[14'd2964] <= 32'h3cd99725;
        mem[14'd2965] <= 32'h3e120274;
        mem[14'd2966] <= 32'h3e2aea0e;
        mem[14'd2967] <= 32'h3e08011a;
        mem[14'd2968] <= 32'h3ef3179b;
        mem[14'd2969] <= 32'h3f21078e;
        mem[14'd2970] <= 32'h3e22a73f;
        mem[14'd2971] <= 32'h3bcc2c2e;
        mem[14'd2972] <= 32'hbc8fb181;
        mem[14'd2973] <= 32'h3c412e0b;
        mem[14'd2974] <= 32'h3c0f5b56;
        mem[14'd2975] <= 32'h3dc00e7a;
        mem[14'd2976] <= 32'h3eb9b748;
        mem[14'd2977] <= 32'h3ec9f329;
        mem[14'd2978] <= 32'h3e618f5d;
        mem[14'd2979] <= 32'h3eb1b098;
        mem[14'd2980] <= 32'h3df38bd9;
        mem[14'd2981] <= 32'h3db850de;
        mem[14'd2982] <= 32'h3e7a8cf7;
        mem[14'd2983] <= 32'h3e08e8c7;
        mem[14'd2984] <= 32'h3ea09c07;
        mem[14'd2985] <= 32'h3e768697;
        mem[14'd2986] <= 32'h3dfc8f0f;
        mem[14'd2987] <= 32'hbd22a8c1;
        mem[14'd2988] <= 32'h3dbf5061;
        mem[14'd2989] <= 32'h3e3d92cf;
        mem[14'd2990] <= 32'h3dc104c5;
        mem[14'd2991] <= 32'h3d8306e2;
        mem[14'd2992] <= 32'hbc31ffd8;
        mem[14'd2993] <= 32'h3e01791e;
        mem[14'd2994] <= 32'h3e45a2f0;
        mem[14'd2995] <= 32'h3ec8aae1;
        mem[14'd2996] <= 32'h3f19a6cc;
        mem[14'd2997] <= 32'h3ee1f3c1;
        mem[14'd2998] <= 32'h3d5fe08f;
        mem[14'd2999] <= 32'h3ca0bfe7;
        mem[14'd3000] <= 32'hbc1747aa;
        mem[14'd3001] <= 32'hbba40f24;
        mem[14'd3002] <= 32'hbb9c0f54;
        mem[14'd3003] <= 32'h3af2f534;
        mem[14'd3004] <= 32'h3e81d8ca;
        mem[14'd3005] <= 32'h3e5401b8;
        mem[14'd3006] <= 32'h3e225126;
        mem[14'd3007] <= 32'h3ead2a91;
        mem[14'd3008] <= 32'h3e72525f;
        mem[14'd3009] <= 32'h3e79b42c;
        mem[14'd3010] <= 32'h3e837c58;
        mem[14'd3011] <= 32'h3e68b987;
        mem[14'd3012] <= 32'h3e5fe9cd;
        mem[14'd3013] <= 32'h3e97ea72;
        mem[14'd3014] <= 32'h3e04f1c5;
        mem[14'd3015] <= 32'h3deafff3;
        mem[14'd3016] <= 32'h3e1b37c5;
        mem[14'd3017] <= 32'h3e2f2080;
        mem[14'd3018] <= 32'h3d8b50a1;
        mem[14'd3019] <= 32'hbc756d72;
        mem[14'd3020] <= 32'h3dcb302e;
        mem[14'd3021] <= 32'h3e523d28;
        mem[14'd3022] <= 32'h3e9e2cf7;
        mem[14'd3023] <= 32'h3e9a4c55;
        mem[14'd3024] <= 32'h3ea07f7d;
        mem[14'd3025] <= 32'h3e9d082a;
        mem[14'd3026] <= 32'h3dc13e00;
        mem[14'd3027] <= 32'h3c45f9c6;
        mem[14'd3028] <= 32'h3c329e9d;
        mem[14'd3029] <= 32'h3c3e399d;
        mem[14'd3030] <= 32'hba4bebdd;
        mem[14'd3031] <= 32'h3d60e5eb;
        mem[14'd3032] <= 32'h3e83f9e6;
        mem[14'd3033] <= 32'h3e664c1a;
        mem[14'd3034] <= 32'h3e6c2c8a;
        mem[14'd3035] <= 32'h3ec1bc70;
        mem[14'd3036] <= 32'h3e80c867;
        mem[14'd3037] <= 32'h3e7224c7;
        mem[14'd3038] <= 32'h3e52c56a;
        mem[14'd3039] <= 32'h3e994d6f;
        mem[14'd3040] <= 32'h3e22e680;
        mem[14'd3041] <= 32'h3dba089f;
        mem[14'd3042] <= 32'h3ccbaac4;
        mem[14'd3043] <= 32'h3d81c1b2;
        mem[14'd3044] <= 32'h3d90206c;
        mem[14'd3045] <= 32'hbd328efc;
        mem[14'd3046] <= 32'h3df7e31b;
        mem[14'd3047] <= 32'h3e69297e;
        mem[14'd3048] <= 32'h3e505360;
        mem[14'd3049] <= 32'h3e8d7723;
        mem[14'd3050] <= 32'h3e853e42;
        mem[14'd3051] <= 32'h3e980cc9;
        mem[14'd3052] <= 32'h3ea34357;
        mem[14'd3053] <= 32'h3e1311fc;
        mem[14'd3054] <= 32'h3d11af95;
        mem[14'd3055] <= 32'hbc5c2407;
        mem[14'd3056] <= 32'hbac50c54;
        mem[14'd3057] <= 32'hbbf1e3c6;
        mem[14'd3058] <= 32'h3d13db40;
        mem[14'd3059] <= 32'h3da265a6;
        mem[14'd3060] <= 32'h3e0ec2b0;
        mem[14'd3061] <= 32'h3e39791c;
        mem[14'd3062] <= 32'h3e379e87;
        mem[14'd3063] <= 32'h3e150299;
        mem[14'd3064] <= 32'h3d2162ec;
        mem[14'd3065] <= 32'h3e7029bd;
        mem[14'd3066] <= 32'h3e098dee;
        mem[14'd3067] <= 32'h3e07b2c6;
        mem[14'd3068] <= 32'h3d899a6a;
        mem[14'd3069] <= 32'h3db1529f;
        mem[14'd3070] <= 32'h3d06d865;
        mem[14'd3071] <= 32'hbd7d0089;
        mem[14'd3072] <= 32'h3db06ae4;
        mem[14'd3073] <= 32'h3e2c7f9e;
        mem[14'd3074] <= 32'h3e856fc1;
        mem[14'd3075] <= 32'h3eaaa129;
        mem[14'd3076] <= 32'h3dd3a9d7;
        mem[14'd3077] <= 32'h3e3e459e;
        mem[14'd3078] <= 32'h3e965f33;
        mem[14'd3079] <= 32'h3ec2dc16;
        mem[14'd3080] <= 32'h3e6afa32;
        mem[14'd3081] <= 32'h3dc62bc5;
        mem[14'd3082] <= 32'h384f2b54;
        mem[14'd3083] <= 32'h3c052b5c;
        mem[14'd3084] <= 32'h3bec437e;
        mem[14'd3085] <= 32'h3bbe94f2;
        mem[14'd3086] <= 32'h3cab67cb;
        mem[14'd3087] <= 32'h3d587157;
        mem[14'd3088] <= 32'h3dea9563;
        mem[14'd3089] <= 32'h3dff0895;
        mem[14'd3090] <= 32'h3e5eb0b7;
        mem[14'd3091] <= 32'h3e7e32e7;
        mem[14'd3092] <= 32'h3e9665bc;
        mem[14'd3093] <= 32'h3e853a3e;
        mem[14'd3094] <= 32'h3e0facec;
        mem[14'd3095] <= 32'h3e036a4c;
        mem[14'd3096] <= 32'h3daa99f0;
        mem[14'd3097] <= 32'hbcc58f25;
        mem[14'd3098] <= 32'hbd6156d7;
        mem[14'd3099] <= 32'hbe048660;
        mem[14'd3100] <= 32'hbcb68393;
        mem[14'd3101] <= 32'h3c979226;
        mem[14'd3102] <= 32'h3e48af46;
        mem[14'd3103] <= 32'h3e492ae6;
        mem[14'd3104] <= 32'h3e778725;
        mem[14'd3105] <= 32'h3e79fa39;
        mem[14'd3106] <= 32'h3e9ae6a8;
        mem[14'd3107] <= 32'h3e5e6c02;
        mem[14'd3108] <= 32'h3e02b0cf;
        mem[14'd3109] <= 32'h3d2f6b71;
        mem[14'd3110] <= 32'hbc07af13;
        mem[14'd3111] <= 32'hba973b30;
        mem[14'd3112] <= 32'hbb536dde;
        mem[14'd3113] <= 32'hbbb1d2fb;
        mem[14'd3114] <= 32'h3c087826;
        mem[14'd3115] <= 32'hbca4d20c;
        mem[14'd3116] <= 32'h3b6d5b76;
        mem[14'd3117] <= 32'hbd4b1a7c;
        mem[14'd3118] <= 32'hbc211e68;
        mem[14'd3119] <= 32'h3d9f94f7;
        mem[14'd3120] <= 32'h3dcadfdb;
        mem[14'd3121] <= 32'h3da56ff8;
        mem[14'd3122] <= 32'h3c853900;
        mem[14'd3123] <= 32'h3dc0ca37;
        mem[14'd3124] <= 32'h3d8ee74f;
        mem[14'd3125] <= 32'hbd47c6cc;
        mem[14'd3126] <= 32'hbd0d9da1;
        mem[14'd3127] <= 32'hbd86944b;
        mem[14'd3128] <= 32'hbd8720eb;
        mem[14'd3129] <= 32'hbcf21bab;
        mem[14'd3130] <= 32'h3e51f3d6;
        mem[14'd3131] <= 32'h3e9c302d;
        mem[14'd3132] <= 32'h3e782229;
        mem[14'd3133] <= 32'h3e8c72aa;
        mem[14'd3134] <= 32'h3e7727f4;
        mem[14'd3135] <= 32'h3e23c190;
        mem[14'd3136] <= 32'h3dcd6ca8;
        mem[14'd3137] <= 32'h3d42e449;
        mem[14'd3138] <= 32'hbc53ecb1;
        mem[14'd3139] <= 32'hba9ef67c;
        mem[14'd3140] <= 32'hbadf66c4;
        mem[14'd3141] <= 32'hbba791fc;
        mem[14'd3142] <= 32'hbaefc152;
        mem[14'd3143] <= 32'hbd2193aa;
        mem[14'd3144] <= 32'hbd7b51c1;
        mem[14'd3145] <= 32'hbe270f97;
        mem[14'd3146] <= 32'hbe80a300;
        mem[14'd3147] <= 32'hbe6bd007;
        mem[14'd3148] <= 32'hbe339663;
        mem[14'd3149] <= 32'hbe156c7b;
        mem[14'd3150] <= 32'hbe53124d;
        mem[14'd3151] <= 32'hbe0c7e5c;
        mem[14'd3152] <= 32'hbc4ddf06;
        mem[14'd3153] <= 32'hbb8a8740;
        mem[14'd3154] <= 32'h3dfbcdb6;
        mem[14'd3155] <= 32'h3c992635;
        mem[14'd3156] <= 32'hbc39524b;
        mem[14'd3157] <= 32'h3dc815af;
        mem[14'd3158] <= 32'h3e013f10;
        mem[14'd3159] <= 32'h3c84c769;
        mem[14'd3160] <= 32'h3cadcc7f;
        mem[14'd3161] <= 32'h3dafd1aa;
        mem[14'd3162] <= 32'h3d11e292;
        mem[14'd3163] <= 32'h3d1cd09d;
        mem[14'd3164] <= 32'h3dc3f41a;
        mem[14'd3165] <= 32'h3d35ba8b;
        mem[14'd3166] <= 32'h3c0dd581;
        mem[14'd3167] <= 32'hbbec9cbd;
        mem[14'd3168] <= 32'h3ba3cd9e;
        mem[14'd3169] <= 32'hbc5d4452;
        mem[14'd3170] <= 32'h3b498ad7;
        mem[14'd3171] <= 32'h3b61078e;
        mem[14'd3172] <= 32'hbcdafa44;
        mem[14'd3173] <= 32'hbd66bb56;
        mem[14'd3174] <= 32'hbd9f54c3;
        mem[14'd3175] <= 32'hbdf7b230;
        mem[14'd3176] <= 32'hbe6c8416;
        mem[14'd3177] <= 32'hbe813cc1;
        mem[14'd3178] <= 32'hbe666d82;
        mem[14'd3179] <= 32'hbe67133b;
        mem[14'd3180] <= 32'hbe15bf4e;
        mem[14'd3181] <= 32'hbe032306;
        mem[14'd3182] <= 32'hbd834eb2;
        mem[14'd3183] <= 32'hbd07fb4f;
        mem[14'd3184] <= 32'hbd7c1e83;
        mem[14'd3185] <= 32'hbd924cc1;
        mem[14'd3186] <= 32'hbddc218e;
        mem[14'd3187] <= 32'hbdfe68f6;
        mem[14'd3188] <= 32'hbdb4fddc;
        mem[14'd3189] <= 32'hbdb72650;
        mem[14'd3190] <= 32'hbd2faa6f;
        mem[14'd3191] <= 32'hbd21b3fd;
        mem[14'd3192] <= 32'hbbdb41c7;
        mem[14'd3193] <= 32'h3ba0b45f;
        mem[14'd3194] <= 32'h3c7e12d0;
        mem[14'd3195] <= 32'hbc8074dc;
        mem[14'd3196] <= 32'hbbc2bc01;
        mem[14'd3197] <= 32'hbc302cfd;
        mem[14'd3198] <= 32'hbc2efc96;
        mem[14'd3199] <= 32'h3c106b24;
        mem[14'd3200] <= 32'h3bbe0512;
        mem[14'd3201] <= 32'hbb85aa59;
        mem[14'd3202] <= 32'hbc91eb2e;
        mem[14'd3203] <= 32'hbcdd6be1;
        mem[14'd3204] <= 32'hbc2240d4;
        mem[14'd3205] <= 32'hbc8a95df;
        mem[14'd3206] <= 32'hbccc8047;
        mem[14'd3207] <= 32'hbcdcaa7f;
        mem[14'd3208] <= 32'hbd1818d6;
        mem[14'd3209] <= 32'hbd3393a2;
        mem[14'd3210] <= 32'hbd09ace0;
        mem[14'd3211] <= 32'hbd64aeec;
        mem[14'd3212] <= 32'hbd7022f7;
        mem[14'd3213] <= 32'hbd295088;
        mem[14'd3214] <= 32'hbd06d71c;
        mem[14'd3215] <= 32'hbc4db928;
        mem[14'd3216] <= 32'hbd03f903;
        mem[14'd3217] <= 32'hbc9361ce;
        mem[14'd3218] <= 32'hbbe66b7f;
        mem[14'd3219] <= 32'hbb0986a5;
        mem[14'd3220] <= 32'h39322577;
        mem[14'd3221] <= 32'hbc137aa8;
        mem[14'd3222] <= 32'h3a24d33a;
        mem[14'd3223] <= 32'h3befd3ec;
        mem[14'd3224] <= 32'h3bf03098;
        mem[14'd3225] <= 32'h3b345ddb;
        mem[14'd3226] <= 32'hbc1cbf2b;
        mem[14'd3227] <= 32'hbca430a1;
        mem[14'd3228] <= 32'hbae3d166;
        mem[14'd3229] <= 32'hbba27751;
        mem[14'd3230] <= 32'hbb95e0fe;
        mem[14'd3231] <= 32'h3b3154c2;
        mem[14'd3232] <= 32'h3c25cd12;
        mem[14'd3233] <= 32'hbc99511d;
        mem[14'd3234] <= 32'h3bc82fb4;
        mem[14'd3235] <= 32'h3c20c680;
        mem[14'd3236] <= 32'hbb124110;
        mem[14'd3237] <= 32'h3bd546f4;
        mem[14'd3238] <= 32'hbbdddcf6;
        mem[14'd3239] <= 32'hbb5ea31d;
        mem[14'd3240] <= 32'h3cadc7cd;
        mem[14'd3241] <= 32'hbba8aaab;
        mem[14'd3242] <= 32'h3ba009a4;
        mem[14'd3243] <= 32'hbcafab8a;
        mem[14'd3244] <= 32'hbca224ba;
        mem[14'd3245] <= 32'h3bc46101;
        mem[14'd3246] <= 32'hbadef180;
        mem[14'd3247] <= 32'h3b3bdbde;
        mem[14'd3248] <= 32'hbbb4ad72;
        mem[14'd3249] <= 32'h3c13f5b0;
        mem[14'd3250] <= 32'hbc5eba7c;
        mem[14'd3251] <= 32'hbb48e07e;
        mem[14'd3252] <= 32'h3b697f9b;
        mem[14'd3253] <= 32'hbb464c69;
        mem[14'd3254] <= 32'hbc1702b0;
        mem[14'd3255] <= 32'hbb974fa6;
        mem[14'd3256] <= 32'h3bb10938;
        mem[14'd3257] <= 32'hbbd62c34;
        mem[14'd3258] <= 32'hba24f5c2;
        mem[14'd3259] <= 32'hbb42b445;
        mem[14'd3260] <= 32'hbc241565;
        mem[14'd3261] <= 32'h3c64f800;
        mem[14'd3262] <= 32'hbae1a984;
        mem[14'd3263] <= 32'h3c6cf7b0;
        mem[14'd3264] <= 32'hbb7afc42;
        mem[14'd3265] <= 32'hbb4063c3;
        mem[14'd3266] <= 32'hbabffc97;
        mem[14'd3267] <= 32'h3c21097a;
        mem[14'd3268] <= 32'hbc1ce67d;
        mem[14'd3269] <= 32'h3a5c7e0f;
        mem[14'd3270] <= 32'h3a87349e;
        mem[14'd3271] <= 32'hb986675f;
        mem[14'd3272] <= 32'hbb605d10;
        mem[14'd3273] <= 32'hbbf35286;
        mem[14'd3274] <= 32'h3c50423d;
        mem[14'd3275] <= 32'hbcb8041d;
        mem[14'd3276] <= 32'h3c161438;
        mem[14'd3277] <= 32'hbc235bc2;
        mem[14'd3278] <= 32'h3bccdaa0;
        mem[14'd3279] <= 32'hbc017b89;
        mem[14'd3280] <= 32'h3c11781b;
        mem[14'd3281] <= 32'hbb580f39;
        mem[14'd3282] <= 32'h3c7f8a25;
        mem[14'd3283] <= 32'hbc8ad924;
        mem[14'd3284] <= 32'hbad2cab2;
        mem[14'd3285] <= 32'hbc053271;
        mem[14'd3286] <= 32'hb916befb;
        mem[14'd3287] <= 32'h3c1d71de;
        mem[14'd3288] <= 32'h3a9f8e74;
        mem[14'd3289] <= 32'hbc503256;
        mem[14'd3290] <= 32'hbc2735ad;
        mem[14'd3291] <= 32'h3c11dba2;
        mem[14'd3292] <= 32'hbbff54ec;
        mem[14'd3293] <= 32'hbc4244b0;
        mem[14'd3294] <= 32'hbbb58491;
        mem[14'd3295] <= 32'hbb8c511e;
        mem[14'd3296] <= 32'hbb292a8e;
        mem[14'd3297] <= 32'h3bd3f4c7;
        mem[14'd3298] <= 32'h3c3ba714;
        mem[14'd3299] <= 32'hbb855813;
        mem[14'd3300] <= 32'hbadac17f;
        mem[14'd3301] <= 32'h3b9e2db2;
        mem[14'd3302] <= 32'h3c144a3a;
        mem[14'd3303] <= 32'h39e27db9;
        mem[14'd3304] <= 32'h3c7830be;
        mem[14'd3305] <= 32'h3bb764a6;
        mem[14'd3306] <= 32'h3bc8d495;
        mem[14'd3307] <= 32'h3cc708d5;
        mem[14'd3308] <= 32'h3b878b4f;
        mem[14'd3309] <= 32'hbc0fc8de;
        mem[14'd3310] <= 32'h3c562cc0;
        mem[14'd3311] <= 32'hbc2ca3c1;
        mem[14'd3312] <= 32'hbb80beb9;
        mem[14'd3313] <= 32'h3c517d07;
        mem[14'd3314] <= 32'hbc37fa39;
        mem[14'd3315] <= 32'hba0b7376;
        mem[14'd3316] <= 32'hbbdec64d;
        mem[14'd3317] <= 32'hbc6d45b6;
        mem[14'd3318] <= 32'hbc8b1d81;
        mem[14'd3319] <= 32'h3abb130d;
        mem[14'd3320] <= 32'h3bfa955a;
        mem[14'd3321] <= 32'h3c0773b0;
        mem[14'd3322] <= 32'hbc9a51a4;
        mem[14'd3323] <= 32'hbc56617a;
        mem[14'd3324] <= 32'hbc322882;
        mem[14'd3325] <= 32'hbcae27fa;
        mem[14'd3326] <= 32'hbced1524;
        mem[14'd3327] <= 32'hbc10ead2;
        mem[14'd3328] <= 32'h3c884ae5;
        mem[14'd3329] <= 32'h3c191124;
        mem[14'd3330] <= 32'h3c4b36fa;
        mem[14'd3331] <= 32'h3b0e873c;
        mem[14'd3332] <= 32'hbb78e72f;
        mem[14'd3333] <= 32'h3c020276;
        mem[14'd3334] <= 32'h3bb147d8;
        mem[14'd3335] <= 32'hbb1609b2;
        mem[14'd3336] <= 32'h3c86c0ec;
        mem[14'd3337] <= 32'hbca1fec9;
        mem[14'd3338] <= 32'h3bf27916;
        mem[14'd3339] <= 32'h3bf68143;
        mem[14'd3340] <= 32'h3a686223;
        mem[14'd3341] <= 32'h3cef10de;
        mem[14'd3342] <= 32'h3cde4fa5;
        mem[14'd3343] <= 32'h3d4f5d1d;
        mem[14'd3344] <= 32'h3d55b416;
        mem[14'd3345] <= 32'h3c6802a3;
        mem[14'd3346] <= 32'h3d81add2;
        mem[14'd3347] <= 32'h3e506514;
        mem[14'd3348] <= 32'h3e91aafb;
        mem[14'd3349] <= 32'h3e6bd4f9;
        mem[14'd3350] <= 32'h3e9854af;
        mem[14'd3351] <= 32'h3e8e5195;
        mem[14'd3352] <= 32'h3e710565;
        mem[14'd3353] <= 32'h3e737825;
        mem[14'd3354] <= 32'h3e49aa60;
        mem[14'd3355] <= 32'h3e07bb1f;
        mem[14'd3356] <= 32'h3ddcf5e1;
        mem[14'd3357] <= 32'hbd0f6cba;
        mem[14'd3358] <= 32'hbd6edf75;
        mem[14'd3359] <= 32'hbcdd2cf7;
        mem[14'd3360] <= 32'hbbc2a12e;
        mem[14'd3361] <= 32'h3ba99288;
        mem[14'd3362] <= 32'hbcb47008;
        mem[14'd3363] <= 32'hbadfd2bc;
        mem[14'd3364] <= 32'h3bf43dd7;
        mem[14'd3365] <= 32'hbc0d72df;
        mem[14'd3366] <= 32'hba2e65f0;
        mem[14'd3367] <= 32'h3b8e7de9;
        mem[14'd3368] <= 32'h3d1f2fc1;
        mem[14'd3369] <= 32'h3dfcee3a;
        mem[14'd3370] <= 32'h3e31f71c;
        mem[14'd3371] <= 32'h3e64ffc0;
        mem[14'd3372] <= 32'h3e987181;
        mem[14'd3373] <= 32'h3e8b3e18;
        mem[14'd3374] <= 32'h3eb2578b;
        mem[14'd3375] <= 32'h3ec82f85;
        mem[14'd3376] <= 32'h3ec48cf0;
        mem[14'd3377] <= 32'h3ec7ef30;
        mem[14'd3378] <= 32'h3e95550f;
        mem[14'd3379] <= 32'h3e950f7f;
        mem[14'd3380] <= 32'h3e9de209;
        mem[14'd3381] <= 32'h3e362d37;
        mem[14'd3382] <= 32'h3e81a0b7;
        mem[14'd3383] <= 32'h3df89622;
        mem[14'd3384] <= 32'hbc99eba6;
        mem[14'd3385] <= 32'hbdecfd20;
        mem[14'd3386] <= 32'hbdfe4c95;
        mem[14'd3387] <= 32'hbe0c9880;
        mem[14'd3388] <= 32'hbcfc3d3a;
        mem[14'd3389] <= 32'hbbd2ee92;
        mem[14'd3390] <= 32'hbc64cbf2;
        mem[14'd3391] <= 32'h3bde42b5;
        mem[14'd3392] <= 32'h3c2d7f84;
        mem[14'd3393] <= 32'hbbedaeec;
        mem[14'd3394] <= 32'h3b109b15;
        mem[14'd3395] <= 32'h3d1c47c7;
        mem[14'd3396] <= 32'h3e04d9de;
        mem[14'd3397] <= 32'h3e832a44;
        mem[14'd3398] <= 32'h3ea006d2;
        mem[14'd3399] <= 32'h3e88e3df;
        mem[14'd3400] <= 32'h3e425c4d;
        mem[14'd3401] <= 32'h3e46339b;
        mem[14'd3402] <= 32'h3e47894a;
        mem[14'd3403] <= 32'h3e286ece;
        mem[14'd3404] <= 32'h3dcce86f;
        mem[14'd3405] <= 32'h3dc4a814;
        mem[14'd3406] <= 32'h3d19de25;
        mem[14'd3407] <= 32'h3e151743;
        mem[14'd3408] <= 32'h3e6bc3c4;
        mem[14'd3409] <= 32'hbcbc625d;
        mem[14'd3410] <= 32'h3cc24fa4;
        mem[14'd3411] <= 32'h3d33d820;
        mem[14'd3412] <= 32'hbda15eda;
        mem[14'd3413] <= 32'hbe39b482;
        mem[14'd3414] <= 32'hbe355a80;
        mem[14'd3415] <= 32'hbe4b7121;
        mem[14'd3416] <= 32'hbd9f3ee7;
        mem[14'd3417] <= 32'hbbf2dd9f;
        mem[14'd3418] <= 32'h3c2bb55d;
        mem[14'd3419] <= 32'h3c4e8587;
        mem[14'd3420] <= 32'h3c4e92de;
        mem[14'd3421] <= 32'hbbd28ecf;
        mem[14'd3422] <= 32'h3c2d3592;
        mem[14'd3423] <= 32'h3dad87dd;
        mem[14'd3424] <= 32'h3e270617;
        mem[14'd3425] <= 32'h3e6e98c1;
        mem[14'd3426] <= 32'h3e8d7f44;
        mem[14'd3427] <= 32'h3e1f0a8c;
        mem[14'd3428] <= 32'h3e030e72;
        mem[14'd3429] <= 32'h3e74fbb7;
        mem[14'd3430] <= 32'h3e83e469;
        mem[14'd3431] <= 32'h3dec00b4;
        mem[14'd3432] <= 32'h3d9337f0;
        mem[14'd3433] <= 32'h3e7a5df1;
        mem[14'd3434] <= 32'h3ddd45b9;
        mem[14'd3435] <= 32'h3e0e63ad;
        mem[14'd3436] <= 32'h3e56b257;
        mem[14'd3437] <= 32'h3d80933d;
        mem[14'd3438] <= 32'h3e38162b;
        mem[14'd3439] <= 32'hbd3064fa;
        mem[14'd3440] <= 32'h3d2b196c;
        mem[14'd3441] <= 32'hbc9963b0;
        mem[14'd3442] <= 32'hbe09dead;
        mem[14'd3443] <= 32'hbe36075a;
        mem[14'd3444] <= 32'hbdf93fd6;
        mem[14'd3445] <= 32'hbd2961d2;
        mem[14'd3446] <= 32'h3bd3e01d;
        mem[14'd3447] <= 32'h3a439572;
        mem[14'd3448] <= 32'h3c22b84d;
        mem[14'd3449] <= 32'h3c26b911;
        mem[14'd3450] <= 32'hbc1f60b2;
        mem[14'd3451] <= 32'h3d83f17c;
        mem[14'd3452] <= 32'h3e86bb89;
        mem[14'd3453] <= 32'h3e95d1ef;
        mem[14'd3454] <= 32'h3e4d6588;
        mem[14'd3455] <= 32'h3d950bb0;
        mem[14'd3456] <= 32'h3d7d5ab7;
        mem[14'd3457] <= 32'h3da8555a;
        mem[14'd3458] <= 32'h3c2e7d98;
        mem[14'd3459] <= 32'hbb0a4258;
        mem[14'd3460] <= 32'h3e0e03a8;
        mem[14'd3461] <= 32'h3d933bea;
        mem[14'd3462] <= 32'h3e71d1ec;
        mem[14'd3463] <= 32'h3e5fd7c8;
        mem[14'd3464] <= 32'h3d14dde4;
        mem[14'd3465] <= 32'h3e0c771a;
        mem[14'd3466] <= 32'h3d18ac2d;
        mem[14'd3467] <= 32'h3dc25e02;
        mem[14'd3468] <= 32'h3d44a15c;
        mem[14'd3469] <= 32'hbddc0f6d;
        mem[14'd3470] <= 32'hbe0713a5;
        mem[14'd3471] <= 32'hbe6ab255;
        mem[14'd3472] <= 32'hbe2f44b2;
        mem[14'd3473] <= 32'hbd2a6abf;
        mem[14'd3474] <= 32'hbc509f74;
        mem[14'd3475] <= 32'h3a9c8d40;
        mem[14'd3476] <= 32'hbc8fc236;
        mem[14'd3477] <= 32'h3bdb6abb;
        mem[14'd3478] <= 32'hbbcf306f;
        mem[14'd3479] <= 32'h3d865f4a;
        mem[14'd3480] <= 32'h3e9f925e;
        mem[14'd3481] <= 32'h3e805c1d;
        mem[14'd3482] <= 32'h3def43e0;
        mem[14'd3483] <= 32'h3d8c6d92;
        mem[14'd3484] <= 32'hbc6022ea;
        mem[14'd3485] <= 32'hbcd2f615;
        mem[14'd3486] <= 32'h3d8ccb5c;
        mem[14'd3487] <= 32'h3ca58abe;
        mem[14'd3488] <= 32'h3dffbb27;
        mem[14'd3489] <= 32'h3dde6dfa;
        mem[14'd3490] <= 32'h3e42611d;
        mem[14'd3491] <= 32'h3e40a911;
        mem[14'd3492] <= 32'h3df001db;
        mem[14'd3493] <= 32'h3def2143;
        mem[14'd3494] <= 32'h3e6975d5;
        mem[14'd3495] <= 32'h3df058b3;
        mem[14'd3496] <= 32'h3dfe121c;
        mem[14'd3497] <= 32'h3dba86b1;
        mem[14'd3498] <= 32'h3de41a4e;
        mem[14'd3499] <= 32'hbe9d6a81;
        mem[14'd3500] <= 32'hbe829bf4;
        mem[14'd3501] <= 32'hbd58e657;
        mem[14'd3502] <= 32'hba6bc8a2;
        mem[14'd3503] <= 32'hbcd62fd7;
        mem[14'd3504] <= 32'hbc50633d;
        mem[14'd3505] <= 32'hbc7a824c;
        mem[14'd3506] <= 32'h3b333a48;
        mem[14'd3507] <= 32'h3dfdf89c;
        mem[14'd3508] <= 32'h3e9f5317;
        mem[14'd3509] <= 32'h3e29d3a5;
        mem[14'd3510] <= 32'h3e18ac06;
        mem[14'd3511] <= 32'h3e02fa0d;
        mem[14'd3512] <= 32'h3d949756;
        mem[14'd3513] <= 32'hbc8c5eca;
        mem[14'd3514] <= 32'hbde81912;
        mem[14'd3515] <= 32'hbea58163;
        mem[14'd3516] <= 32'hbe5f58e3;
        mem[14'd3517] <= 32'hbda21da6;
        mem[14'd3518] <= 32'h3e6b9730;
        mem[14'd3519] <= 32'h3eba4fee;
        mem[14'd3520] <= 32'h3e86e4a6;
        mem[14'd3521] <= 32'h3e1abc30;
        mem[14'd3522] <= 32'h3ddf302a;
        mem[14'd3523] <= 32'h3e23632d;
        mem[14'd3524] <= 32'h3e841aed;
        mem[14'd3525] <= 32'h3e566b73;
        mem[14'd3526] <= 32'h3e478730;
        mem[14'd3527] <= 32'hbe2cb55b;
        mem[14'd3528] <= 32'hbe738e8e;
        mem[14'd3529] <= 32'hbd4d0cee;
        mem[14'd3530] <= 32'hbc6b8143;
        mem[14'd3531] <= 32'h3761576c;
        mem[14'd3532] <= 32'h3aa6410f;
        mem[14'd3533] <= 32'h3c102b41;
        mem[14'd3534] <= 32'h3bf103be;
        mem[14'd3535] <= 32'h3e14e74b;
        mem[14'd3536] <= 32'h3e0b06c9;
        mem[14'd3537] <= 32'hbc2f73a0;
        mem[14'd3538] <= 32'hbccddf86;
        mem[14'd3539] <= 32'hbdbef70f;
        mem[14'd3540] <= 32'hbe73b4a1;
        mem[14'd3541] <= 32'hbed45b58;
        mem[14'd3542] <= 32'hbeecfb3e;
        mem[14'd3543] <= 32'hbef48fd2;
        mem[14'd3544] <= 32'hbedada9e;
        mem[14'd3545] <= 32'h3c04543e;
        mem[14'd3546] <= 32'h3e3fa899;
        mem[14'd3547] <= 32'h3e434a04;
        mem[14'd3548] <= 32'h3e6e1430;
        mem[14'd3549] <= 32'h3e3ba0bd;
        mem[14'd3550] <= 32'h3e2b484c;
        mem[14'd3551] <= 32'h3e574836;
        mem[14'd3552] <= 32'h3e86422e;
        mem[14'd3553] <= 32'h3e1ea6a3;
        mem[14'd3554] <= 32'h3da282a2;
        mem[14'd3555] <= 32'hbdbdc3ee;
        mem[14'd3556] <= 32'hbe1ec393;
        mem[14'd3557] <= 32'hbd1c875a;
        mem[14'd3558] <= 32'hbc4f7821;
        mem[14'd3559] <= 32'hbb550691;
        mem[14'd3560] <= 32'h3c59f84e;
        mem[14'd3561] <= 32'hbbb70072;
        mem[14'd3562] <= 32'h3cbfd4cd;
        mem[14'd3563] <= 32'h3de6abbc;
        mem[14'd3564] <= 32'h3d6e829c;
        mem[14'd3565] <= 32'hbe24aa1a;
        mem[14'd3566] <= 32'hbe8272c9;
        mem[14'd3567] <= 32'hbed1d0e1;
        mem[14'd3568] <= 32'hbeee62b9;
        mem[14'd3569] <= 32'hbedb896a;
        mem[14'd3570] <= 32'hbea6f5ba;
        mem[14'd3571] <= 32'hbe3b4db4;
        mem[14'd3572] <= 32'hbdb05696;
        mem[14'd3573] <= 32'h3df99c81;
        mem[14'd3574] <= 32'h3e55e910;
        mem[14'd3575] <= 32'h3e3e7c2b;
        mem[14'd3576] <= 32'h3ca6a6ff;
        mem[14'd3577] <= 32'h3e753085;
        mem[14'd3578] <= 32'h3def78b9;
        mem[14'd3579] <= 32'h3e27b4f5;
        mem[14'd3580] <= 32'h3e81df6d;
        mem[14'd3581] <= 32'hbd3c2110;
        mem[14'd3582] <= 32'hbd91a713;
        mem[14'd3583] <= 32'hbe0751a6;
        mem[14'd3584] <= 32'hbdfc6b5c;
        mem[14'd3585] <= 32'hbb5b406e;
        mem[14'd3586] <= 32'hbcb935af;
        mem[14'd3587] <= 32'hbcb8ac44;
        mem[14'd3588] <= 32'hbc826376;
        mem[14'd3589] <= 32'h3a841be1;
        mem[14'd3590] <= 32'hbc4838b1;
        mem[14'd3591] <= 32'h3cd143af;
        mem[14'd3592] <= 32'hbd710593;
        mem[14'd3593] <= 32'hbe5851dd;
        mem[14'd3594] <= 32'hbeadabf4;
        mem[14'd3595] <= 32'hbeb3e6a8;
        mem[14'd3596] <= 32'hbeaeb9a8;
        mem[14'd3597] <= 32'hbe0c0170;
        mem[14'd3598] <= 32'h3d6c570e;
        mem[14'd3599] <= 32'hbd7bfafd;
        mem[14'd3600] <= 32'h3d7b96aa;
        mem[14'd3601] <= 32'h3e03d1b9;
        mem[14'd3602] <= 32'h3eb8c3b0;
        mem[14'd3603] <= 32'h3e1624f2;
        mem[14'd3604] <= 32'h3dc467d8;
        mem[14'd3605] <= 32'h3d97cbf3;
        mem[14'd3606] <= 32'h3e1b2c7d;
        mem[14'd3607] <= 32'h3c932596;
        mem[14'd3608] <= 32'hbdd5012b;
        mem[14'd3609] <= 32'hbeb300df;
        mem[14'd3610] <= 32'hbe95ac62;
        mem[14'd3611] <= 32'hbe176871;
        mem[14'd3612] <= 32'hbd923fa7;
        mem[14'd3613] <= 32'hbb17539e;
        mem[14'd3614] <= 32'hbb8ef71b;
        mem[14'd3615] <= 32'h3b900f73;
        mem[14'd3616] <= 32'hba3cb08a;
        mem[14'd3617] <= 32'hbc3a1a59;
        mem[14'd3618] <= 32'hbcbb1db4;
        mem[14'd3619] <= 32'hbc14939b;
        mem[14'd3620] <= 32'hbdfc4c8f;
        mem[14'd3621] <= 32'hbe748476;
        mem[14'd3622] <= 32'hbe9b67ac;
        mem[14'd3623] <= 32'hbe9d02c4;
        mem[14'd3624] <= 32'hbe3e6f02;
        mem[14'd3625] <= 32'hbdaec37e;
        mem[14'd3626] <= 32'hbe14c9e7;
        mem[14'd3627] <= 32'hbe4846c0;
        mem[14'd3628] <= 32'h3d909137;
        mem[14'd3629] <= 32'h3e9686ae;
        mem[14'd3630] <= 32'h3e73f095;
        mem[14'd3631] <= 32'hbda84fc3;
        mem[14'd3632] <= 32'h3d6dde67;
        mem[14'd3633] <= 32'h3db7b5d3;
        mem[14'd3634] <= 32'h3e28c7f2;
        mem[14'd3635] <= 32'hbdb84042;
        mem[14'd3636] <= 32'hbea9ac81;
        mem[14'd3637] <= 32'hbeb6e25d;
        mem[14'd3638] <= 32'hbeb68c6c;
        mem[14'd3639] <= 32'hbe3c8380;
        mem[14'd3640] <= 32'hbd5a1839;
        mem[14'd3641] <= 32'hbc8abae7;
        mem[14'd3642] <= 32'h3b4bdf11;
        mem[14'd3643] <= 32'hbc3684e1;
        mem[14'd3644] <= 32'h3c11047e;
        mem[14'd3645] <= 32'hba8785c6;
        mem[14'd3646] <= 32'h3bd0944d;
        mem[14'd3647] <= 32'h39af46e8;
        mem[14'd3648] <= 32'hbd7678fa;
        mem[14'd3649] <= 32'hbe67db6c;
        mem[14'd3650] <= 32'hbe9dc712;
        mem[14'd3651] <= 32'hbeafe2c3;
        mem[14'd3652] <= 32'hbe46228f;
        mem[14'd3653] <= 32'hbd885d71;
        mem[14'd3654] <= 32'hbe12a271;
        mem[14'd3655] <= 32'hbe386987;
        mem[14'd3656] <= 32'h3db6b972;
        mem[14'd3657] <= 32'h3dc08f3a;
        mem[14'd3658] <= 32'h3dcf17e4;
        mem[14'd3659] <= 32'h3d21fbcd;
        mem[14'd3660] <= 32'hbcb9124c;
        mem[14'd3661] <= 32'h3d2fc885;
        mem[14'd3662] <= 32'h3d12af3d;
        mem[14'd3663] <= 32'hbdb88d34;
        mem[14'd3664] <= 32'hbe251f73;
        mem[14'd3665] <= 32'hbd9284ba;
        mem[14'd3666] <= 32'hbe5979a4;
        mem[14'd3667] <= 32'hbde942c9;
        mem[14'd3668] <= 32'hbd6a6c4c;
        mem[14'd3669] <= 32'hbc92738f;
        mem[14'd3670] <= 32'h3c1e3e37;
        mem[14'd3671] <= 32'h3c01775d;
        mem[14'd3672] <= 32'hbc9a9bef;
        mem[14'd3673] <= 32'h3cdfdfa6;
        mem[14'd3674] <= 32'h3d144cda;
        mem[14'd3675] <= 32'h3b6023b0;
        mem[14'd3676] <= 32'h3b9b4950;
        mem[14'd3677] <= 32'hbd9d5dd1;
        mem[14'd3678] <= 32'hbe27c62d;
        mem[14'd3679] <= 32'hbe88f8d4;
        mem[14'd3680] <= 32'hbe8f712f;
        mem[14'd3681] <= 32'hbe592026;
        mem[14'd3682] <= 32'hbe351440;
        mem[14'd3683] <= 32'hbd86b2bc;
        mem[14'd3684] <= 32'h3d52e689;
        mem[14'd3685] <= 32'h3df6d303;
        mem[14'd3686] <= 32'h3e165b17;
        mem[14'd3687] <= 32'h3dc7a48d;
        mem[14'd3688] <= 32'hbcd92e3e;
        mem[14'd3689] <= 32'hbd15ffc3;
        mem[14'd3690] <= 32'hbda1d6ae;
        mem[14'd3691] <= 32'h3db84aff;
        mem[14'd3692] <= 32'h3e4e8c1d;
        mem[14'd3693] <= 32'h3e1b6d60;
        mem[14'd3694] <= 32'h3e1dc2f7;
        mem[14'd3695] <= 32'h3dfb7343;
        mem[14'd3696] <= 32'h3d2dc80e;
        mem[14'd3697] <= 32'hbd5f869c;
        mem[14'd3698] <= 32'h3bfc0b00;
        mem[14'd3699] <= 32'hbad2c40e;
        mem[14'd3700] <= 32'hbbe415c9;
        mem[14'd3701] <= 32'h3cc12724;
        mem[14'd3702] <= 32'h3d4a8a1f;
        mem[14'd3703] <= 32'h3da91d3f;
        mem[14'd3704] <= 32'h3e3e2d2d;
        mem[14'd3705] <= 32'h3d460e9a;
        mem[14'd3706] <= 32'hbdd091bc;
        mem[14'd3707] <= 32'hbe62fd5b;
        mem[14'd3708] <= 32'hbeb437ce;
        mem[14'd3709] <= 32'hbe4f01ed;
        mem[14'd3710] <= 32'hbe4a85ac;
        mem[14'd3711] <= 32'hbdb37387;
        mem[14'd3712] <= 32'h3c88897c;
        mem[14'd3713] <= 32'h3e58e499;
        mem[14'd3714] <= 32'hbc0ff23f;
        mem[14'd3715] <= 32'hbe3a8295;
        mem[14'd3716] <= 32'hbe7527b0;
        mem[14'd3717] <= 32'hbd393e75;
        mem[14'd3718] <= 32'h3e488774;
        mem[14'd3719] <= 32'h3e879854;
        mem[14'd3720] <= 32'h3e1d76d8;
        mem[14'd3721] <= 32'h3e1ab043;
        mem[14'd3722] <= 32'h3e7b2fae;
        mem[14'd3723] <= 32'h3e7e631d;
        mem[14'd3724] <= 32'h3df02b6b;
        mem[14'd3725] <= 32'hbd6c3737;
        mem[14'd3726] <= 32'hbb0432ca;
        mem[14'd3727] <= 32'h3b8e6bd9;
        mem[14'd3728] <= 32'hbc49e818;
        mem[14'd3729] <= 32'h3ba2d02c;
        mem[14'd3730] <= 32'h3d5217c2;
        mem[14'd3731] <= 32'h3e4c70f6;
        mem[14'd3732] <= 32'h3e87534a;
        mem[14'd3733] <= 32'h3db6537b;
        mem[14'd3734] <= 32'hbd62d13d;
        mem[14'd3735] <= 32'hbdc1be0c;
        mem[14'd3736] <= 32'hbe69a117;
        mem[14'd3737] <= 32'hbee7cd5e;
        mem[14'd3738] <= 32'hbf04530d;
        mem[14'd3739] <= 32'hbee23e5c;
        mem[14'd3740] <= 32'hbe899849;
        mem[14'd3741] <= 32'hbe574678;
        mem[14'd3742] <= 32'hbeb3d989;
        mem[14'd3743] <= 32'hbe7e310e;
        mem[14'd3744] <= 32'h3cbfb8fb;
        mem[14'd3745] <= 32'h3e3dc581;
        mem[14'd3746] <= 32'h3dc5bd5c;
        mem[14'd3747] <= 32'h3ea6ce27;
        mem[14'd3748] <= 32'h3d26408f;
        mem[14'd3749] <= 32'h3e40dd60;
        mem[14'd3750] <= 32'h3e9721ae;
        mem[14'd3751] <= 32'h3e825c21;
        mem[14'd3752] <= 32'hbd0c67db;
        mem[14'd3753] <= 32'hbdbbb9ad;
        mem[14'd3754] <= 32'h3a9578c3;
        mem[14'd3755] <= 32'h3c5bab52;
        mem[14'd3756] <= 32'h3a6f16f1;
        mem[14'd3757] <= 32'hbc16fd31;
        mem[14'd3758] <= 32'h3d4616a9;
        mem[14'd3759] <= 32'h3eae75a1;
        mem[14'd3760] <= 32'h3ea3c2d9;
        mem[14'd3761] <= 32'h3e8532ec;
        mem[14'd3762] <= 32'h3dce6a75;
        mem[14'd3763] <= 32'hbde7a8f0;
        mem[14'd3764] <= 32'hbdf1fa87;
        mem[14'd3765] <= 32'hbeae743d;
        mem[14'd3766] <= 32'hbed36ae5;
        mem[14'd3767] <= 32'hbec0226a;
        mem[14'd3768] <= 32'hbee5c2f4;
        mem[14'd3769] <= 32'hbeb09a17;
        mem[14'd3770] <= 32'hbe8d7155;
        mem[14'd3771] <= 32'h3dc56d52;
        mem[14'd3772] <= 32'h3e994167;
        mem[14'd3773] <= 32'h3e5db307;
        mem[14'd3774] <= 32'h3e383eda;
        mem[14'd3775] <= 32'h3e591958;
        mem[14'd3776] <= 32'h3dd87534;
        mem[14'd3777] <= 32'h3ea12802;
        mem[14'd3778] <= 32'h3ea86519;
        mem[14'd3779] <= 32'h3ddde90e;
        mem[14'd3780] <= 32'hbe0c5698;
        mem[14'd3781] <= 32'hbd60a547;
        mem[14'd3782] <= 32'h3c8ae900;
        mem[14'd3783] <= 32'h3c92eddf;
        mem[14'd3784] <= 32'hbccb2072;
        mem[14'd3785] <= 32'hbb9effd8;
        mem[14'd3786] <= 32'h3c61db09;
        mem[14'd3787] <= 32'h3eb19703;
        mem[14'd3788] <= 32'h3eb62a92;
        mem[14'd3789] <= 32'h3ecb3681;
        mem[14'd3790] <= 32'h3e2e62e3;
        mem[14'd3791] <= 32'h3cf09135;
        mem[14'd3792] <= 32'h3b99a916;
        mem[14'd3793] <= 32'hbd1cc11c;
        mem[14'd3794] <= 32'hbdfbb8d0;
        mem[14'd3795] <= 32'hbe6898a3;
        mem[14'd3796] <= 32'hbe745357;
        mem[14'd3797] <= 32'hbe189973;
        mem[14'd3798] <= 32'hbd2eb24a;
        mem[14'd3799] <= 32'h3d9e9e99;
        mem[14'd3800] <= 32'h3e1f888c;
        mem[14'd3801] <= 32'h3e8d2442;
        mem[14'd3802] <= 32'h3e60a995;
        mem[14'd3803] <= 32'h3e37146d;
        mem[14'd3804] <= 32'h3d941e36;
        mem[14'd3805] <= 32'h3e907618;
        mem[14'd3806] <= 32'h3e23f28a;
        mem[14'd3807] <= 32'h3d1ce01e;
        mem[14'd3808] <= 32'hbdbfbbc5;
        mem[14'd3809] <= 32'hbd605c39;
        mem[14'd3810] <= 32'hbb5bda63;
        mem[14'd3811] <= 32'h3ba1c76d;
        mem[14'd3812] <= 32'h38575abd;
        mem[14'd3813] <= 32'hbb8fd291;
        mem[14'd3814] <= 32'h3ccc589d;
        mem[14'd3815] <= 32'h3e9f1cdf;
        mem[14'd3816] <= 32'h3eb3a739;
        mem[14'd3817] <= 32'h3e966e33;
        mem[14'd3818] <= 32'h3ea02104;
        mem[14'd3819] <= 32'h3e3eeb05;
        mem[14'd3820] <= 32'h3e38a93e;
        mem[14'd3821] <= 32'h3e4d233f;
        mem[14'd3822] <= 32'hbd017182;
        mem[14'd3823] <= 32'hbe3a936c;
        mem[14'd3824] <= 32'hbea20314;
        mem[14'd3825] <= 32'hbdd99501;
        mem[14'd3826] <= 32'h3d2bc21d;
        mem[14'd3827] <= 32'hbc66b8b3;
        mem[14'd3828] <= 32'h3dda11d4;
        mem[14'd3829] <= 32'h3e2fd09a;
        mem[14'd3830] <= 32'h3e787433;
        mem[14'd3831] <= 32'h3e03ed6e;
        mem[14'd3832] <= 32'h3e82daa6;
        mem[14'd3833] <= 32'h3df8c9b9;
        mem[14'd3834] <= 32'h3ca08838;
        mem[14'd3835] <= 32'h39e3f3b8;
        mem[14'd3836] <= 32'hbdaab850;
        mem[14'd3837] <= 32'hbca57bc3;
        mem[14'd3838] <= 32'hbbf8a8af;
        mem[14'd3839] <= 32'h3c458d82;
        mem[14'd3840] <= 32'h3bff2b61;
        mem[14'd3841] <= 32'hbb270598;
        mem[14'd3842] <= 32'h3d413d09;
        mem[14'd3843] <= 32'h3e43fcd1;
        mem[14'd3844] <= 32'h3e7b7cfd;
        mem[14'd3845] <= 32'h3dccc6fe;
        mem[14'd3846] <= 32'h3e3f20ae;
        mem[14'd3847] <= 32'h3e13c53f;
        mem[14'd3848] <= 32'h3dd9cd4f;
        mem[14'd3849] <= 32'hbe00e14e;
        mem[14'd3850] <= 32'hbe041880;
        mem[14'd3851] <= 32'hbe074361;
        mem[14'd3852] <= 32'hbdb7dec0;
        mem[14'd3853] <= 32'hbdbb9200;
        mem[14'd3854] <= 32'hbd6f0c91;
        mem[14'd3855] <= 32'hbaca1a7e;
        mem[14'd3856] <= 32'h3dde7fb7;
        mem[14'd3857] <= 32'h3d82428f;
        mem[14'd3858] <= 32'h3e422a2d;
        mem[14'd3859] <= 32'h3e7dc5c7;
        mem[14'd3860] <= 32'h3d830335;
        mem[14'd3861] <= 32'hbd4a317b;
        mem[14'd3862] <= 32'hbd54a4c0;
        mem[14'd3863] <= 32'hbe033cd4;
        mem[14'd3864] <= 32'hbdf4d4b4;
        mem[14'd3865] <= 32'hbcf23899;
        mem[14'd3866] <= 32'hbb3b57fc;
        mem[14'd3867] <= 32'hbc5eff86;
        mem[14'd3868] <= 32'hbc4e7266;
        mem[14'd3869] <= 32'hb91ad1aa;
        mem[14'd3870] <= 32'h3d41be99;
        mem[14'd3871] <= 32'h3e04f8cc;
        mem[14'd3872] <= 32'h3e3a11eb;
        mem[14'd3873] <= 32'h3e014010;
        mem[14'd3874] <= 32'h3dbf971c;
        mem[14'd3875] <= 32'h3d173eca;
        mem[14'd3876] <= 32'hbd199f57;
        mem[14'd3877] <= 32'h3c4e85e8;
        mem[14'd3878] <= 32'h3c4a59a2;
        mem[14'd3879] <= 32'h3db45b60;
        mem[14'd3880] <= 32'hbda4abd3;
        mem[14'd3881] <= 32'hbda4b76d;
        mem[14'd3882] <= 32'hbdac74e0;
        mem[14'd3883] <= 32'h3d865ac5;
        mem[14'd3884] <= 32'h3cfab1e4;
        mem[14'd3885] <= 32'h3dcc5cbd;
        mem[14'd3886] <= 32'h3db085fe;
        mem[14'd3887] <= 32'h3e23ccfd;
        mem[14'd3888] <= 32'h3d937df0;
        mem[14'd3889] <= 32'hbd8727ac;
        mem[14'd3890] <= 32'hbcfc09e2;
        mem[14'd3891] <= 32'hbd8923eb;
        mem[14'd3892] <= 32'hbd71647e;
        mem[14'd3893] <= 32'hbc01b525;
        mem[14'd3894] <= 32'hbc3478fb;
        mem[14'd3895] <= 32'hbc53c4c0;
        mem[14'd3896] <= 32'h3ca88e66;
        mem[14'd3897] <= 32'hbb74cb72;
        mem[14'd3898] <= 32'h3cfcda2d;
        mem[14'd3899] <= 32'h3e0b66eb;
        mem[14'd3900] <= 32'h3e6ec1a5;
        mem[14'd3901] <= 32'h3e745c15;
        mem[14'd3902] <= 32'h3e7e8126;
        mem[14'd3903] <= 32'h3e4955c2;
        mem[14'd3904] <= 32'hbb025923;
        mem[14'd3905] <= 32'h3da2d1a0;
        mem[14'd3906] <= 32'h3dd98fb8;
        mem[14'd3907] <= 32'h3de0e0da;
        mem[14'd3908] <= 32'hbdf69984;
        mem[14'd3909] <= 32'h3d5319d7;
        mem[14'd3910] <= 32'hbd84b0cc;
        mem[14'd3911] <= 32'hbd48acad;
        mem[14'd3912] <= 32'hbe05f314;
        mem[14'd3913] <= 32'h3d46a46b;
        mem[14'd3914] <= 32'h3e598bcb;
        mem[14'd3915] <= 32'h3d6382df;
        mem[14'd3916] <= 32'hbd0e67e0;
        mem[14'd3917] <= 32'hbda091bc;
        mem[14'd3918] <= 32'hbdc2bc0f;
        mem[14'd3919] <= 32'hbd88c28b;
        mem[14'd3920] <= 32'hbcc5e881;
        mem[14'd3921] <= 32'hbcc880c4;
        mem[14'd3922] <= 32'hbb27c36d;
        mem[14'd3923] <= 32'h3bf4b3db;
        mem[14'd3924] <= 32'h3a98a514;
        mem[14'd3925] <= 32'h3c920b93;
        mem[14'd3926] <= 32'h3bf87f5e;
        mem[14'd3927] <= 32'h3dbb3744;
        mem[14'd3928] <= 32'h3e50d2cd;
        mem[14'd3929] <= 32'h3e6e4618;
        mem[14'd3930] <= 32'h3eb3f40f;
        mem[14'd3931] <= 32'h3ecd10f4;
        mem[14'd3932] <= 32'h3e994d33;
        mem[14'd3933] <= 32'h3e63b03f;
        mem[14'd3934] <= 32'h3ea3b4ca;
        mem[14'd3935] <= 32'h3e953901;
        mem[14'd3936] <= 32'h3e63b9b6;
        mem[14'd3937] <= 32'h3e9a3811;
        mem[14'd3938] <= 32'h3e716359;
        mem[14'd3939] <= 32'h3df9b79e;
        mem[14'd3940] <= 32'h3e31ec07;
        mem[14'd3941] <= 32'h3dda8c24;
        mem[14'd3942] <= 32'hbd96c63b;
        mem[14'd3943] <= 32'hbdf1cd7a;
        mem[14'd3944] <= 32'hbd874473;
        mem[14'd3945] <= 32'hbccdcb3b;
        mem[14'd3946] <= 32'hbcb7b803;
        mem[14'd3947] <= 32'hbcac5489;
        mem[14'd3948] <= 32'hbc920548;
        mem[14'd3949] <= 32'hbbf1eb30;
        mem[14'd3950] <= 32'hbc57e7d0;
        mem[14'd3951] <= 32'hbc480ee6;
        mem[14'd3952] <= 32'hba9c2e63;
        mem[14'd3953] <= 32'hbc180e14;
        mem[14'd3954] <= 32'h3c7242af;
        mem[14'd3955] <= 32'h39715f9d;
        mem[14'd3956] <= 32'h3cd40e73;
        mem[14'd3957] <= 32'h3d5a81c9;
        mem[14'd3958] <= 32'h3e291833;
        mem[14'd3959] <= 32'h3e8a533c;
        mem[14'd3960] <= 32'h3ed484f3;
        mem[14'd3961] <= 32'h3eed0c05;
        mem[14'd3962] <= 32'h3f01ad46;
        mem[14'd3963] <= 32'h3ee9f985;
        mem[14'd3964] <= 32'h3f012d5d;
        mem[14'd3965] <= 32'h3eda19b3;
        mem[14'd3966] <= 32'h3e868f47;
        mem[14'd3967] <= 32'h3dfd5c69;
        mem[14'd3968] <= 32'h3dfbbbfc;
        mem[14'd3969] <= 32'h3ce8f7ce;
        mem[14'd3970] <= 32'h3d01dad4;
        mem[14'd3971] <= 32'h3d4f2315;
        mem[14'd3972] <= 32'hbc856ec0;
        mem[14'd3973] <= 32'hbcc69499;
        mem[14'd3974] <= 32'hbc15afec;
        mem[14'd3975] <= 32'hbc338569;
        mem[14'd3976] <= 32'h3b63257d;
        mem[14'd3977] <= 32'hbc0ac930;
        mem[14'd3978] <= 32'hbc82e4b6;
        mem[14'd3979] <= 32'hbb597ad5;
        mem[14'd3980] <= 32'h3b77bddb;
        mem[14'd3981] <= 32'h3ad6095b;
        mem[14'd3982] <= 32'hbc37984d;
        mem[14'd3983] <= 32'hbae687aa;
        mem[14'd3984] <= 32'hbc13a207;
        mem[14'd3985] <= 32'h3b4592d0;
        mem[14'd3986] <= 32'hba51c9ba;
        mem[14'd3987] <= 32'h3c492fd8;
        mem[14'd3988] <= 32'hbb112ce1;
        mem[14'd3989] <= 32'h3b2b23df;
        mem[14'd3990] <= 32'h3c6d6af7;
        mem[14'd3991] <= 32'h3c11d22e;
        mem[14'd3992] <= 32'h3ba4bf14;
        mem[14'd3993] <= 32'h3aea8418;
        mem[14'd3994] <= 32'h3bf26cfd;
        mem[14'd3995] <= 32'hbc9fe42f;
        mem[14'd3996] <= 32'h3d06822d;
        mem[14'd3997] <= 32'h3c8644f6;
        mem[14'd3998] <= 32'h3b779c72;
        mem[14'd3999] <= 32'hbbd4cacb;
        mem[14'd4000] <= 32'h3c129d24;
        mem[14'd4001] <= 32'hbc559fad;
        mem[14'd4002] <= 32'hbbabbdf6;
        mem[14'd4003] <= 32'h3aa95a6f;
        mem[14'd4004] <= 32'h3c8696b6;
        mem[14'd4005] <= 32'h3c05dd30;
        mem[14'd4006] <= 32'h3c111a8a;
        mem[14'd4007] <= 32'hbc87e6f1;
        mem[14'd4008] <= 32'hbb2914a1;
        mem[14'd4009] <= 32'hbbf29b77;
        mem[14'd4010] <= 32'h3c23797b;
        mem[14'd4011] <= 32'h3c74e0dc;
        mem[14'd4012] <= 32'hbbd9d164;
        mem[14'd4013] <= 32'h3b658180;
        mem[14'd4014] <= 32'h3c61b21e;
        mem[14'd4015] <= 32'h3bb8532c;
        mem[14'd4016] <= 32'hbbb4846d;
        mem[14'd4017] <= 32'hbc862f75;
        mem[14'd4018] <= 32'hbbabad41;
        mem[14'd4019] <= 32'hbbd7f477;
        mem[14'd4020] <= 32'hbcc8012c;
        mem[14'd4021] <= 32'h3aaf727f;
        mem[14'd4022] <= 32'hbbdc4c51;
        mem[14'd4023] <= 32'hbbb73f18;
        mem[14'd4024] <= 32'h3c34c8ed;
        mem[14'd4025] <= 32'hbba6c1df;
        mem[14'd4026] <= 32'hbbe96373;
        mem[14'd4027] <= 32'hbcf90b36;
        mem[14'd4028] <= 32'hbb498a22;
        mem[14'd4029] <= 32'h3c0cd2dc;
        mem[14'd4030] <= 32'h3ba8ec58;
        mem[14'd4031] <= 32'h3b9bde8f;
        mem[14'd4032] <= 32'h3ca3ed80;
        mem[14'd4033] <= 32'h3c64f1e1;
        mem[14'd4034] <= 32'hbb8e2533;
        mem[14'd4035] <= 32'hbbf5fa81;
        mem[14'd4036] <= 32'hbcc79f38;
        mem[14'd4037] <= 32'h3c35fe34;
        mem[14'd4038] <= 32'hbcd0082e;
        mem[14'd4039] <= 32'hbac3baa9;
        mem[14'd4040] <= 32'hba493df9;
        mem[14'd4041] <= 32'hbc497ac2;
        mem[14'd4042] <= 32'hbbe23ef0;
        mem[14'd4043] <= 32'hbc6eb6c3;
        mem[14'd4044] <= 32'h3a30a064;
        mem[14'd4045] <= 32'hbbcc24bb;
        mem[14'd4046] <= 32'hbbe2dfaa;
        mem[14'd4047] <= 32'hbb2039eb;
        mem[14'd4048] <= 32'hbc221daa;
        mem[14'd4049] <= 32'hbcbfc4ba;
        mem[14'd4050] <= 32'h38a8003f;
        mem[14'd4051] <= 32'h3ba4dcf2;
        mem[14'd4052] <= 32'hba9fd8d2;
        mem[14'd4053] <= 32'hbc421cfd;
        mem[14'd4054] <= 32'hbbb4a87e;
        mem[14'd4055] <= 32'hbb6f0afc;
        mem[14'd4056] <= 32'h3b25058a;
        mem[14'd4057] <= 32'h3b93cbc8;
        mem[14'd4058] <= 32'hbb56bb93;
        mem[14'd4059] <= 32'h3b6e2b3d;
        mem[14'd4060] <= 32'h3c5141f4;
        mem[14'd4061] <= 32'hbcce94e6;
        mem[14'd4062] <= 32'hbc2a566e;
        mem[14'd4063] <= 32'hbb34c066;
        mem[14'd4064] <= 32'hbc9be469;
        mem[14'd4065] <= 32'hbb100fdb;
        mem[14'd4066] <= 32'hbc31bc65;
        mem[14'd4067] <= 32'h3b280e85;
        mem[14'd4068] <= 32'hbb926306;
        mem[14'd4069] <= 32'h3bb20630;
        mem[14'd4070] <= 32'hbc8697fc;
        mem[14'd4071] <= 32'hbd360cd8;
        mem[14'd4072] <= 32'hbd23704b;
        mem[14'd4073] <= 32'hbc9e9da6;
        mem[14'd4074] <= 32'hbd0e7874;
        mem[14'd4075] <= 32'hbd2abc0a;
        mem[14'd4076] <= 32'hbdaf30bc;
        mem[14'd4077] <= 32'hbd56cac8;
        mem[14'd4078] <= 32'hbcacb2de;
        mem[14'd4079] <= 32'hbd80c1da;
        mem[14'd4080] <= 32'hbd8b4ae6;
        mem[14'd4081] <= 32'hbd0482ab;
        mem[14'd4082] <= 32'hbc8fe080;
        mem[14'd4083] <= 32'hbd162575;
        mem[14'd4084] <= 32'hbd04375a;
        mem[14'd4085] <= 32'hbcc3288f;
        mem[14'd4086] <= 32'hbc84b636;
        mem[14'd4087] <= 32'hbbf1430d;
        mem[14'd4088] <= 32'hbb31f2c2;
        mem[14'd4089] <= 32'h3b3e25c7;
        mem[14'd4090] <= 32'hbb396e15;
        mem[14'd4091] <= 32'hb94a9d38;
        mem[14'd4092] <= 32'hbc7fed29;
        mem[14'd4093] <= 32'hbc968480;
        mem[14'd4094] <= 32'hbba84c36;
        mem[14'd4095] <= 32'hbca82655;
        mem[14'd4096] <= 32'hbc9f0301;
        mem[14'd4097] <= 32'h3c2eaf65;
        mem[14'd4098] <= 32'hbd01de96;
        mem[14'd4099] <= 32'hbd40aea1;
        mem[14'd4100] <= 32'hbd9630ee;
        mem[14'd4101] <= 32'hbd8a8b9e;
        mem[14'd4102] <= 32'hbe11a093;
        mem[14'd4103] <= 32'hbe1eed84;
        mem[14'd4104] <= 32'hbe549159;
        mem[14'd4105] <= 32'hbe3fd8af;
        mem[14'd4106] <= 32'hbe04f1f6;
        mem[14'd4107] <= 32'hbe0fe01d;
        mem[14'd4108] <= 32'hbe1f523f;
        mem[14'd4109] <= 32'hbdac1325;
        mem[14'd4110] <= 32'hbd668338;
        mem[14'd4111] <= 32'hbd549bf9;
        mem[14'd4112] <= 32'hbd0331f5;
        mem[14'd4113] <= 32'hbcb6dbf0;
        mem[14'd4114] <= 32'hbd180546;
        mem[14'd4115] <= 32'hbc2b0308;
        mem[14'd4116] <= 32'hbbc14848;
        mem[14'd4117] <= 32'h3c561d40;
        mem[14'd4118] <= 32'hbbacb710;
        mem[14'd4119] <= 32'h3bb9b601;
        mem[14'd4120] <= 32'hbbb97490;
        mem[14'd4121] <= 32'h3ae7237b;
        mem[14'd4122] <= 32'hbc2c603f;
        mem[14'd4123] <= 32'hbbf1aa72;
        mem[14'd4124] <= 32'h3acfc368;
        mem[14'd4125] <= 32'hbbb1957d;
        mem[14'd4126] <= 32'hbca8b812;
        mem[14'd4127] <= 32'hbd86d803;
        mem[14'd4128] <= 32'hbdeb8bc9;
        mem[14'd4129] <= 32'hbe38f804;
        mem[14'd4130] <= 32'hbe73e9ca;
        mem[14'd4131] <= 32'hbe947b03;
        mem[14'd4132] <= 32'hbeb80f0c;
        mem[14'd4133] <= 32'hbedbfbeb;
        mem[14'd4134] <= 32'hbeb98249;
        mem[14'd4135] <= 32'hbeb7d84c;
        mem[14'd4136] <= 32'hbe90a850;
        mem[14'd4137] <= 32'hbe56de04;
        mem[14'd4138] <= 32'hbe0d02dc;
        mem[14'd4139] <= 32'hbd0e836c;
        mem[14'd4140] <= 32'hbb1eaeb8;
        mem[14'd4141] <= 32'h3c920721;
        mem[14'd4142] <= 32'h3b704d04;
        mem[14'd4143] <= 32'h3c3fbd60;
        mem[14'd4144] <= 32'h3b8a7e48;
        mem[14'd4145] <= 32'hbbbe8f27;
        mem[14'd4146] <= 32'h3c5bcfa9;
        mem[14'd4147] <= 32'h3ba20270;
        mem[14'd4148] <= 32'h39d6368c;
        mem[14'd4149] <= 32'h38d24a4d;
        mem[14'd4150] <= 32'h3c5c1370;
        mem[14'd4151] <= 32'h3b65a812;
        mem[14'd4152] <= 32'h3c8ec72c;
        mem[14'd4153] <= 32'h3c1944aa;
        mem[14'd4154] <= 32'hbd2d0b38;
        mem[14'd4155] <= 32'hbd37873d;
        mem[14'd4156] <= 32'hbe06b068;
        mem[14'd4157] <= 32'hbe4c826f;
        mem[14'd4158] <= 32'hbe907380;
        mem[14'd4159] <= 32'hbe937bc2;
        mem[14'd4160] <= 32'hbe9a591d;
        mem[14'd4161] <= 32'hbe86fdb7;
        mem[14'd4162] <= 32'hbe9ab92b;
        mem[14'd4163] <= 32'hbeaf7033;
        mem[14'd4164] <= 32'hbe479671;
        mem[14'd4165] <= 32'hbe20b7ca;
        mem[14'd4166] <= 32'hbdee533a;
        mem[14'd4167] <= 32'h3d506e00;
        mem[14'd4168] <= 32'h3e1cfa13;
        mem[14'd4169] <= 32'h3e181496;
        mem[14'd4170] <= 32'h3e2b3406;
        mem[14'd4171] <= 32'h3e110633;
        mem[14'd4172] <= 32'h3d9a5587;
        mem[14'd4173] <= 32'h3bff5d1d;
        mem[14'd4174] <= 32'hbb9834ca;
        mem[14'd4175] <= 32'h3c0ebaec;
        mem[14'd4176] <= 32'h3c0668bf;
        mem[14'd4177] <= 32'h3ad826b9;
        mem[14'd4178] <= 32'hbaa8f2da;
        mem[14'd4179] <= 32'hbb8041dd;
        mem[14'd4180] <= 32'h3bad5e63;
        mem[14'd4181] <= 32'h3d6edf41;
        mem[14'd4182] <= 32'h3cf7de6e;
        mem[14'd4183] <= 32'hbc5fadd8;
        mem[14'd4184] <= 32'hbccfa344;
        mem[14'd4185] <= 32'hbd1b446b;
        mem[14'd4186] <= 32'hbdfca9f9;
        mem[14'd4187] <= 32'hbe209d63;
        mem[14'd4188] <= 32'hbe1d3b6f;
        mem[14'd4189] <= 32'hbe7b18e2;
        mem[14'd4190] <= 32'hbda209e6;
        mem[14'd4191] <= 32'hbd85cc08;
        mem[14'd4192] <= 32'h3c69724e;
        mem[14'd4193] <= 32'hbc8bd075;
        mem[14'd4194] <= 32'h3d361dda;
        mem[14'd4195] <= 32'h3dda36a8;
        mem[14'd4196] <= 32'h3dc0a6c1;
        mem[14'd4197] <= 32'h3dc25eeb;
        mem[14'd4198] <= 32'h3e55f58f;
        mem[14'd4199] <= 32'h3e9f5f76;
        mem[14'd4200] <= 32'h3dee97ac;
        mem[14'd4201] <= 32'hbc3d6dc3;
        mem[14'd4202] <= 32'hbc69b0c4;
        mem[14'd4203] <= 32'h3c584998;
        mem[14'd4204] <= 32'hbc178f17;
        mem[14'd4205] <= 32'hbaaefa99;
        mem[14'd4206] <= 32'hbc6a1212;
        mem[14'd4207] <= 32'hbca9ea8d;
        mem[14'd4208] <= 32'h3d0680e9;
        mem[14'd4209] <= 32'h3de3b918;
        mem[14'd4210] <= 32'h3da91e6a;
        mem[14'd4211] <= 32'h3d95e18e;
        mem[14'd4212] <= 32'h3ceb4d75;
        mem[14'd4213] <= 32'h3ca7f4e5;
        mem[14'd4214] <= 32'hbdbd4596;
        mem[14'd4215] <= 32'hbe3e2ec9;
        mem[14'd4216] <= 32'hbe532f0c;
        mem[14'd4217] <= 32'hbe9e2f87;
        mem[14'd4218] <= 32'hbea275ad;
        mem[14'd4219] <= 32'hbeb49e86;
        mem[14'd4220] <= 32'hbe96876d;
        mem[14'd4221] <= 32'hbe553e73;
        mem[14'd4222] <= 32'hbe7c2c86;
        mem[14'd4223] <= 32'hbd6bc18d;
        mem[14'd4224] <= 32'hbd82cc03;
        mem[14'd4225] <= 32'h3c712c65;
        mem[14'd4226] <= 32'h3e8d0f8b;
        mem[14'd4227] <= 32'h3ec0128d;
        mem[14'd4228] <= 32'h3e09d5a4;
        mem[14'd4229] <= 32'h3b528a72;
        mem[14'd4230] <= 32'h3b5fc9cb;
        mem[14'd4231] <= 32'h3c1a7b40;
        mem[14'd4232] <= 32'hbc7ba9f5;
        mem[14'd4233] <= 32'hbbf9ba69;
        mem[14'd4234] <= 32'hbaf3fb04;
        mem[14'd4235] <= 32'hbbbc2f39;
        mem[14'd4236] <= 32'h3cf6ee3d;
        mem[14'd4237] <= 32'h3e0e8172;
        mem[14'd4238] <= 32'h3d8a42e8;
        mem[14'd4239] <= 32'h3d4c5456;
        mem[14'd4240] <= 32'hbceba56a;
        mem[14'd4241] <= 32'hbcec2c34;
        mem[14'd4242] <= 32'hbe1aeaae;
        mem[14'd4243] <= 32'hbe4dbb30;
        mem[14'd4244] <= 32'hbec450e4;
        mem[14'd4245] <= 32'hbeab07a6;
        mem[14'd4246] <= 32'hbec7a785;
        mem[14'd4247] <= 32'hbeca2938;
        mem[14'd4248] <= 32'hbed01ba7;
        mem[14'd4249] <= 32'hbe613387;
        mem[14'd4250] <= 32'hbe54cdea;
        mem[14'd4251] <= 32'hbdf705a9;
        mem[14'd4252] <= 32'hbe01a584;
        mem[14'd4253] <= 32'hbcc4c4cc;
        mem[14'd4254] <= 32'h3e1b0647;
        mem[14'd4255] <= 32'h3e9ece5e;
        mem[14'd4256] <= 32'h3df6db71;
        mem[14'd4257] <= 32'h3d1a79ec;
        mem[14'd4258] <= 32'h3d36382d;
        mem[14'd4259] <= 32'h3c2c37ec;
        mem[14'd4260] <= 32'hbcb6d2da;
        mem[14'd4261] <= 32'hbb67812b;
        mem[14'd4262] <= 32'hbbe5e59a;
        mem[14'd4263] <= 32'hbc40430b;
        mem[14'd4264] <= 32'h3caba527;
        mem[14'd4265] <= 32'h3dc4f0d5;
        mem[14'd4266] <= 32'h3cec487c;
        mem[14'd4267] <= 32'h3c26339d;
        mem[14'd4268] <= 32'hbde9e8f3;
        mem[14'd4269] <= 32'hbc9f50c6;
        mem[14'd4270] <= 32'hbe1316f1;
        mem[14'd4271] <= 32'hbe0a495c;
        mem[14'd4272] <= 32'hbe81b840;
        mem[14'd4273] <= 32'hbe7ba698;
        mem[14'd4274] <= 32'hbec2df12;
        mem[14'd4275] <= 32'hbebd42e0;
        mem[14'd4276] <= 32'hbeba72fd;
        mem[14'd4277] <= 32'hbe69f00f;
        mem[14'd4278] <= 32'hbdafbe94;
        mem[14'd4279] <= 32'hbd8a1c45;
        mem[14'd4280] <= 32'hbdb24876;
        mem[14'd4281] <= 32'hbd2e241e;
        mem[14'd4282] <= 32'hbc958f51;
        mem[14'd4283] <= 32'h3dd686fe;
        mem[14'd4284] <= 32'h3cea7857;
        mem[14'd4285] <= 32'h3c6dc544;
        mem[14'd4286] <= 32'hbcc1cdaf;
        mem[14'd4287] <= 32'hbb00f145;
        mem[14'd4288] <= 32'h3b1e4e98;
        mem[14'd4289] <= 32'h3ba7686a;
        mem[14'd4290] <= 32'hbbc5d72b;
        mem[14'd4291] <= 32'hbda4e18a;
        mem[14'd4292] <= 32'hbdac3032;
        mem[14'd4293] <= 32'hbc16e270;
        mem[14'd4294] <= 32'hbd9ad54a;
        mem[14'd4295] <= 32'hbdaa3158;
        mem[14'd4296] <= 32'hbd794863;
        mem[14'd4297] <= 32'hbd6ccd80;
        mem[14'd4298] <= 32'hbe1398d4;
        mem[14'd4299] <= 32'hbdc09ec8;
        mem[14'd4300] <= 32'hbdf0d25a;
        mem[14'd4301] <= 32'hbe153cc7;
        mem[14'd4302] <= 32'hbf16e8c3;
        mem[14'd4303] <= 32'hbebcaab5;
        mem[14'd4304] <= 32'hbd9d311d;
        mem[14'd4305] <= 32'hbdbe0a7e;
        mem[14'd4306] <= 32'h3c8e69c0;
        mem[14'd4307] <= 32'h3bb142eb;
        mem[14'd4308] <= 32'hbbd6976e;
        mem[14'd4309] <= 32'hbba488d7;
        mem[14'd4310] <= 32'hbcd7d36a;
        mem[14'd4311] <= 32'hbd98d539;
        mem[14'd4312] <= 32'hbe476686;
        mem[14'd4313] <= 32'hbe0d3941;
        mem[14'd4314] <= 32'hbd4002aa;
        mem[14'd4315] <= 32'hbc7868c4;
        mem[14'd4316] <= 32'hbc304c03;
        mem[14'd4317] <= 32'hbc85c838;
        mem[14'd4318] <= 32'hbd754543;
        mem[14'd4319] <= 32'hbde433e1;
        mem[14'd4320] <= 32'hbde57194;
        mem[14'd4321] <= 32'hbdd3f864;
        mem[14'd4322] <= 32'hbe14219c;
        mem[14'd4323] <= 32'hbd442dd3;
        mem[14'd4324] <= 32'hbce11baa;
        mem[14'd4325] <= 32'h3e02edc1;
        mem[14'd4326] <= 32'h3d63b481;
        mem[14'd4327] <= 32'h3d465501;
        mem[14'd4328] <= 32'h3e3edc2d;
        mem[14'd4329] <= 32'hbe7cf612;
        mem[14'd4330] <= 32'hbf3c5f23;
        mem[14'd4331] <= 32'hbdfdb3e3;
        mem[14'd4332] <= 32'hbd1de8f6;
        mem[14'd4333] <= 32'h3d52c41a;
        mem[14'd4334] <= 32'hbce448fd;
        mem[14'd4335] <= 32'h3d839949;
        mem[14'd4336] <= 32'hbde89242;
        mem[14'd4337] <= 32'hbd917b0c;
        mem[14'd4338] <= 32'hbdb4c4bc;
        mem[14'd4339] <= 32'hbea7baaa;
        mem[14'd4340] <= 32'hbe8bb49c;
        mem[14'd4341] <= 32'hbe28f45a;
        mem[14'd4342] <= 32'hbd792c68;
        mem[14'd4343] <= 32'hbcb6bd06;
        mem[14'd4344] <= 32'hbb535101;
        mem[14'd4345] <= 32'hbcc02845;
        mem[14'd4346] <= 32'hbd902d31;
        mem[14'd4347] <= 32'hbddebeee;
        mem[14'd4348] <= 32'hbe056a4c;
        mem[14'd4349] <= 32'hbdb1ef01;
        mem[14'd4350] <= 32'hbbba5aa4;
        mem[14'd4351] <= 32'h3d333405;
        mem[14'd4352] <= 32'h3e2d238c;
        mem[14'd4353] <= 32'h3ea6aa2a;
        mem[14'd4354] <= 32'h3eb2ddef;
        mem[14'd4355] <= 32'h3e610fee;
        mem[14'd4356] <= 32'h3ec1fac5;
        mem[14'd4357] <= 32'hbef3c8b5;
        mem[14'd4358] <= 32'hbf287c14;
        mem[14'd4359] <= 32'h3dddc6a8;
        mem[14'd4360] <= 32'h3ea75357;
        mem[14'd4361] <= 32'h3df86fea;
        mem[14'd4362] <= 32'hbd30605f;
        mem[14'd4363] <= 32'hbd109f52;
        mem[14'd4364] <= 32'hbe2c6f2b;
        mem[14'd4365] <= 32'hbdf98499;
        mem[14'd4366] <= 32'hbe26da0e;
        mem[14'd4367] <= 32'hbea359b9;
        mem[14'd4368] <= 32'hbe810c86;
        mem[14'd4369] <= 32'hbdec9577;
        mem[14'd4370] <= 32'hbcc64a65;
        mem[14'd4371] <= 32'hbb45b972;
        mem[14'd4372] <= 32'hbb552082;
        mem[14'd4373] <= 32'hbcfa415f;
        mem[14'd4374] <= 32'hbd6245fc;
        mem[14'd4375] <= 32'hbe08e141;
        mem[14'd4376] <= 32'hbe35a9b4;
        mem[14'd4377] <= 32'hbcf2d832;
        mem[14'd4378] <= 32'h3dcbb40a;
        mem[14'd4379] <= 32'h3e9469c6;
        mem[14'd4380] <= 32'h3eb3801c;
        mem[14'd4381] <= 32'h3e960d22;
        mem[14'd4382] <= 32'h3ed66deb;
        mem[14'd4383] <= 32'h3f09d9c0;
        mem[14'd4384] <= 32'h3f296d3b;
        mem[14'd4385] <= 32'hbd89df08;
        mem[14'd4386] <= 32'hbec2ea76;
        mem[14'd4387] <= 32'h3e585903;
        mem[14'd4388] <= 32'h3eb9ba7f;
        mem[14'd4389] <= 32'h3d5410d5;
        mem[14'd4390] <= 32'hbbbce927;
        mem[14'd4391] <= 32'h3da98cd0;
        mem[14'd4392] <= 32'h3d95fd49;
        mem[14'd4393] <= 32'h3e10f992;
        mem[14'd4394] <= 32'h3b3a588c;
        mem[14'd4395] <= 32'hbe1a5002;
        mem[14'd4396] <= 32'hbda62761;
        mem[14'd4397] <= 32'hbd2f8439;
        mem[14'd4398] <= 32'hbc57e7b3;
        mem[14'd4399] <= 32'hbbe525a5;
        mem[14'd4400] <= 32'hbc613b79;
        mem[14'd4401] <= 32'hbcad2fc8;
        mem[14'd4402] <= 32'hbd48bd01;
        mem[14'd4403] <= 32'hbdbd4228;
        mem[14'd4404] <= 32'hbd3d1592;
        mem[14'd4405] <= 32'h3e09c9e2;
        mem[14'd4406] <= 32'h3ea10455;
        mem[14'd4407] <= 32'h3eb48998;
        mem[14'd4408] <= 32'h3ea7b960;
        mem[14'd4409] <= 32'h3ea64fa4;
        mem[14'd4410] <= 32'h3ed44892;
        mem[14'd4411] <= 32'h3f1dd5bc;
        mem[14'd4412] <= 32'h3ed86768;
        mem[14'd4413] <= 32'hbe2a629f;
        mem[14'd4414] <= 32'hbdde7e50;
        mem[14'd4415] <= 32'h3e8f945e;
        mem[14'd4416] <= 32'h3e80fbb8;
        mem[14'd4417] <= 32'h3e90702b;
        mem[14'd4418] <= 32'h3e62476d;
        mem[14'd4419] <= 32'h3e2bdf24;
        mem[14'd4420] <= 32'h3e9b4c9a;
        mem[14'd4421] <= 32'h3e7252de;
        mem[14'd4422] <= 32'h3e0e31f0;
        mem[14'd4423] <= 32'hbd851706;
        mem[14'd4424] <= 32'hbdeaa660;
        mem[14'd4425] <= 32'hbc7d58af;
        mem[14'd4426] <= 32'hbd073b39;
        mem[14'd4427] <= 32'h3c7be7db;
        mem[14'd4428] <= 32'hbacef2c8;
        mem[14'd4429] <= 32'hbc08a7cd;
        mem[14'd4430] <= 32'hbc9ff93a;
        mem[14'd4431] <= 32'hbc6810ca;
        mem[14'd4432] <= 32'h3e54414a;
        mem[14'd4433] <= 32'h3eb106a4;
        mem[14'd4434] <= 32'h3ead66eb;
        mem[14'd4435] <= 32'h3eb0d95d;
        mem[14'd4436] <= 32'h3e9c2d23;
        mem[14'd4437] <= 32'h3e6ea3f7;
        mem[14'd4438] <= 32'h3e8fb488;
        mem[14'd4439] <= 32'h3ecd41b5;
        mem[14'd4440] <= 32'h3e7eda94;
        mem[14'd4441] <= 32'hbe1fd266;
        mem[14'd4442] <= 32'hbd074289;
        mem[14'd4443] <= 32'h3e2b2534;
        mem[14'd4444] <= 32'h3ec63e85;
        mem[14'd4445] <= 32'h3ef2d4fa;
        mem[14'd4446] <= 32'h3e882efd;
        mem[14'd4447] <= 32'h3ec4746e;
        mem[14'd4448] <= 32'h3e3e9d8d;
        mem[14'd4449] <= 32'h3de0d0af;
        mem[14'd4450] <= 32'h3dd71002;
        mem[14'd4451] <= 32'hbd56cb5f;
        mem[14'd4452] <= 32'hbe03516b;
        mem[14'd4453] <= 32'hbd0f0659;
        mem[14'd4454] <= 32'hbd303eb0;
        mem[14'd4455] <= 32'h3a659dbc;
        mem[14'd4456] <= 32'h3bc7e846;
        mem[14'd4457] <= 32'h3b0111c0;
        mem[14'd4458] <= 32'h3b7dcc47;
        mem[14'd4459] <= 32'h3d005d26;
        mem[14'd4460] <= 32'h3e1690a0;
        mem[14'd4461] <= 32'h3e27fa87;
        mem[14'd4462] <= 32'h3e620059;
        mem[14'd4463] <= 32'h3e9d7a05;
        mem[14'd4464] <= 32'h3ea637f6;
        mem[14'd4465] <= 32'h3e9fbd60;
        mem[14'd4466] <= 32'h3e670a52;
        mem[14'd4467] <= 32'h3e9934b3;
        mem[14'd4468] <= 32'h3e146349;
        mem[14'd4469] <= 32'hbe0d0b7e;
        mem[14'd4470] <= 32'h3d06cbc1;
        mem[14'd4471] <= 32'h3e8a557c;
        mem[14'd4472] <= 32'h3efaa4ab;
        mem[14'd4473] <= 32'h3ebe5bab;
        mem[14'd4474] <= 32'h3e110242;
        mem[14'd4475] <= 32'h3e30bff6;
        mem[14'd4476] <= 32'hbd2bf718;
        mem[14'd4477] <= 32'hbcc4086e;
        mem[14'd4478] <= 32'h3d92d6dc;
        mem[14'd4479] <= 32'hbda6ace8;
        mem[14'd4480] <= 32'hbe77be7d;
        mem[14'd4481] <= 32'hbde5a8f7;
        mem[14'd4482] <= 32'hbc91c579;
        mem[14'd4483] <= 32'h3b058802;
        mem[14'd4484] <= 32'hbbe79e53;
        mem[14'd4485] <= 32'hbc0bbf5a;
        mem[14'd4486] <= 32'hbbba16f4;
        mem[14'd4487] <= 32'hbd879fdd;
        mem[14'd4488] <= 32'hbdfdcaf3;
        mem[14'd4489] <= 32'hba36cc46;
        mem[14'd4490] <= 32'h3dd877f1;
        mem[14'd4491] <= 32'h3ea2d680;
        mem[14'd4492] <= 32'h3ebe9eb0;
        mem[14'd4493] <= 32'h3e57e923;
        mem[14'd4494] <= 32'h3c2470e9;
        mem[14'd4495] <= 32'hbd1ac0d2;
        mem[14'd4496] <= 32'h3d3cca58;
        mem[14'd4497] <= 32'h3d35dd59;
        mem[14'd4498] <= 32'h3e865ed0;
        mem[14'd4499] <= 32'h3efee87a;
        mem[14'd4500] <= 32'h3ed58390;
        mem[14'd4501] <= 32'h3ea20a05;
        mem[14'd4502] <= 32'h3e451625;
        mem[14'd4503] <= 32'h3defeab7;
        mem[14'd4504] <= 32'h3e15e5fb;
        mem[14'd4505] <= 32'h3db048b0;
        mem[14'd4506] <= 32'hbd807726;
        mem[14'd4507] <= 32'hbe2186ae;
        mem[14'd4508] <= 32'hbe46fb97;
        mem[14'd4509] <= 32'hbe031605;
        mem[14'd4510] <= 32'hbd734b4a;
        mem[14'd4511] <= 32'h3be0b18d;
        mem[14'd4512] <= 32'hbbbcc659;
        mem[14'd4513] <= 32'hbc8de595;
        mem[14'd4514] <= 32'hbb80a7f9;
        mem[14'd4515] <= 32'hbdfffe5f;
        mem[14'd4516] <= 32'hbe058efc;
        mem[14'd4517] <= 32'hbdd55599;
        mem[14'd4518] <= 32'hbd0e0452;
        mem[14'd4519] <= 32'h3e3c6545;
        mem[14'd4520] <= 32'h3e86c3b2;
        mem[14'd4521] <= 32'h3e03532d;
        mem[14'd4522] <= 32'hbcdda0f3;
        mem[14'd4523] <= 32'hbdb3b137;
        mem[14'd4524] <= 32'h3d3654d8;
        mem[14'd4525] <= 32'h3e8a02e9;
        mem[14'd4526] <= 32'h3ef74834;
        mem[14'd4527] <= 32'h3ec80895;
        mem[14'd4528] <= 32'h3eacafc4;
        mem[14'd4529] <= 32'h3e620e86;
        mem[14'd4530] <= 32'h3e45e7ad;
        mem[14'd4531] <= 32'hbd75ae92;
        mem[14'd4532] <= 32'h3cac4982;
        mem[14'd4533] <= 32'h3d626211;
        mem[14'd4534] <= 32'hbe1d75e4;
        mem[14'd4535] <= 32'hbe0d51bd;
        mem[14'd4536] <= 32'hbe1ec137;
        mem[14'd4537] <= 32'hbe087daa;
        mem[14'd4538] <= 32'hbd3faaad;
        mem[14'd4539] <= 32'hbca6dc75;
        mem[14'd4540] <= 32'h3be6f14d;
        mem[14'd4541] <= 32'hbb03821b;
        mem[14'd4542] <= 32'hbc805f80;
        mem[14'd4543] <= 32'hbdd2dcac;
        mem[14'd4544] <= 32'hbdfc5161;
        mem[14'd4545] <= 32'hbdb083c0;
        mem[14'd4546] <= 32'hbd91a966;
        mem[14'd4547] <= 32'hbba7d7ca;
        mem[14'd4548] <= 32'h3d9403f1;
        mem[14'd4549] <= 32'h3d3386db;
        mem[14'd4550] <= 32'hbe5a4abf;
        mem[14'd4551] <= 32'hbdd5995b;
        mem[14'd4552] <= 32'h3e39d30d;
        mem[14'd4553] <= 32'h3e91926e;
        mem[14'd4554] <= 32'h3e94d1e1;
        mem[14'd4555] <= 32'h3e687b3a;
        mem[14'd4556] <= 32'h3e485455;
        mem[14'd4557] <= 32'hbe0d3cee;
        mem[14'd4558] <= 32'hbdcc9b39;
        mem[14'd4559] <= 32'hbdda18c6;
        mem[14'd4560] <= 32'hbca7afae;
        mem[14'd4561] <= 32'hbda6d08a;
        mem[14'd4562] <= 32'hbe9a028e;
        mem[14'd4563] <= 32'hbe45a31d;
        mem[14'd4564] <= 32'hbe1ab134;
        mem[14'd4565] <= 32'hbdd4a3ee;
        mem[14'd4566] <= 32'h39b8d079;
        mem[14'd4567] <= 32'hba760f89;
        mem[14'd4568] <= 32'hbaaacfa5;
        mem[14'd4569] <= 32'h3a2f060c;
        mem[14'd4570] <= 32'hbcb79275;
        mem[14'd4571] <= 32'hbd1c12fe;
        mem[14'd4572] <= 32'hbdc3fde1;
        mem[14'd4573] <= 32'hbd857316;
        mem[14'd4574] <= 32'hbdc68ea6;
        mem[14'd4575] <= 32'hbe2925a3;
        mem[14'd4576] <= 32'hbe8dcadb;
        mem[14'd4577] <= 32'hbeaa5b68;
        mem[14'd4578] <= 32'hbebdc09e;
        mem[14'd4579] <= 32'hbe620638;
        mem[14'd4580] <= 32'hbea9b6ab;
        mem[14'd4581] <= 32'hbddf2a72;
        mem[14'd4582] <= 32'h3dbbc408;
        mem[14'd4583] <= 32'h3d65ccc7;
        mem[14'd4584] <= 32'hbbe077d6;
        mem[14'd4585] <= 32'hbe08616c;
        mem[14'd4586] <= 32'hbe077da8;
        mem[14'd4587] <= 32'hbe542b12;
        mem[14'd4588] <= 32'hbe273b04;
        mem[14'd4589] <= 32'hbdf6e4c5;
        mem[14'd4590] <= 32'hbe9dc2f4;
        mem[14'd4591] <= 32'hbe7058cd;
        mem[14'd4592] <= 32'hbe0b5213;
        mem[14'd4593] <= 32'hbcfb6d4c;
        mem[14'd4594] <= 32'h3a441311;
        mem[14'd4595] <= 32'hbcd8ea60;
        mem[14'd4596] <= 32'h3c3277c6;
        mem[14'd4597] <= 32'hbbb81b0f;
        mem[14'd4598] <= 32'hbc101baf;
        mem[14'd4599] <= 32'hbd38a636;
        mem[14'd4600] <= 32'hbddfffa4;
        mem[14'd4601] <= 32'hbe2808da;
        mem[14'd4602] <= 32'hbe661fc8;
        mem[14'd4603] <= 32'hbeb407ec;
        mem[14'd4604] <= 32'hbed48fa8;
        mem[14'd4605] <= 32'hbec8e1cc;
        mem[14'd4606] <= 32'hbecb28d7;
        mem[14'd4607] <= 32'hbe584ea1;
        mem[14'd4608] <= 32'hbe6a8b51;
        mem[14'd4609] <= 32'hbeac5cce;
        mem[14'd4610] <= 32'hbdc6d578;
        mem[14'd4611] <= 32'hbc9934e5;
        mem[14'd4612] <= 32'h3c873861;
        mem[14'd4613] <= 32'h3bfb2e46;
        mem[14'd4614] <= 32'hbde878cf;
        mem[14'd4615] <= 32'hbe43b3ce;
        mem[14'd4616] <= 32'hbdf7560c;
        mem[14'd4617] <= 32'hbd8bae97;
        mem[14'd4618] <= 32'hbe309e89;
        mem[14'd4619] <= 32'hbe2ff20b;
        mem[14'd4620] <= 32'hbddc094e;
        mem[14'd4621] <= 32'hbd25987d;
        mem[14'd4622] <= 32'h3c32f7e1;
        mem[14'd4623] <= 32'hbc1396c3;
        mem[14'd4624] <= 32'hbb97e4c0;
        mem[14'd4625] <= 32'h3b0b5920;
        mem[14'd4626] <= 32'h3b9b590d;
        mem[14'd4627] <= 32'hbd23d4fc;
        mem[14'd4628] <= 32'hbdb238a5;
        mem[14'd4629] <= 32'hbdd2b877;
        mem[14'd4630] <= 32'hbe90e8ee;
        mem[14'd4631] <= 32'hbebc6325;
        mem[14'd4632] <= 32'hbe63b37c;
        mem[14'd4633] <= 32'hbe522a0f;
        mem[14'd4634] <= 32'hbe572511;
        mem[14'd4635] <= 32'hbde66bfe;
        mem[14'd4636] <= 32'hbe246119;
        mem[14'd4637] <= 32'hbe5bf289;
        mem[14'd4638] <= 32'hbdf9831e;
        mem[14'd4639] <= 32'hbc94d770;
        mem[14'd4640] <= 32'hbd9ccb82;
        mem[14'd4641] <= 32'h3c8be48f;
        mem[14'd4642] <= 32'hbdbb62c9;
        mem[14'd4643] <= 32'hbbf6fe25;
        mem[14'd4644] <= 32'h3cddd135;
        mem[14'd4645] <= 32'h3c98a3f1;
        mem[14'd4646] <= 32'hbd321b20;
        mem[14'd4647] <= 32'hbda15d2f;
        mem[14'd4648] <= 32'hbd85aed0;
        mem[14'd4649] <= 32'hbd52dea0;
        mem[14'd4650] <= 32'hbacd27d3;
        mem[14'd4651] <= 32'h3b6ce82e;
        mem[14'd4652] <= 32'h3c4d9a15;
        mem[14'd4653] <= 32'hbbf76c2d;
        mem[14'd4654] <= 32'hbc86fee0;
        mem[14'd4655] <= 32'hbd1da67b;
        mem[14'd4656] <= 32'hbd3f6bca;
        mem[14'd4657] <= 32'hbdf08fbd;
        mem[14'd4658] <= 32'hbe22dc8e;
        mem[14'd4659] <= 32'hbe540f71;
        mem[14'd4660] <= 32'hbe491153;
        mem[14'd4661] <= 32'hbe3ecea1;
        mem[14'd4662] <= 32'hbddc9842;
        mem[14'd4663] <= 32'hbdac4376;
        mem[14'd4664] <= 32'hbe1c6a50;
        mem[14'd4665] <= 32'hbdbc6b95;
        mem[14'd4666] <= 32'hbe0e7d38;
        mem[14'd4667] <= 32'hbd947baf;
        mem[14'd4668] <= 32'hbd89b980;
        mem[14'd4669] <= 32'h3d238188;
        mem[14'd4670] <= 32'h3cfb437b;
        mem[14'd4671] <= 32'h3e4ce25d;
        mem[14'd4672] <= 32'h3dffe963;
        mem[14'd4673] <= 32'h3e26db38;
        mem[14'd4674] <= 32'hbb97f7c8;
        mem[14'd4675] <= 32'hbd2a0d35;
        mem[14'd4676] <= 32'hbc9af680;
        mem[14'd4677] <= 32'hbb78c2e7;
        mem[14'd4678] <= 32'hbb94f8fc;
        mem[14'd4679] <= 32'hbb4f07d3;
        mem[14'd4680] <= 32'h3c3225cf;
        mem[14'd4681] <= 32'h3c977db7;
        mem[14'd4682] <= 32'hbc1abc2c;
        mem[14'd4683] <= 32'hbc5db9fe;
        mem[14'd4684] <= 32'hbcba2530;
        mem[14'd4685] <= 32'hbd7927c1;
        mem[14'd4686] <= 32'hbd9c6bdf;
        mem[14'd4687] <= 32'hbda585e4;
        mem[14'd4688] <= 32'hbd52a9e5;
        mem[14'd4689] <= 32'hbbda9e2b;
        mem[14'd4690] <= 32'hbcc30c74;
        mem[14'd4691] <= 32'h3b932995;
        mem[14'd4692] <= 32'hbdbb397d;
        mem[14'd4693] <= 32'hbdabe4ef;
        mem[14'd4694] <= 32'hbd34cb21;
        mem[14'd4695] <= 32'hbcf643d3;
        mem[14'd4696] <= 32'h3d52308e;
        mem[14'd4697] <= 32'h3dadf41d;
        mem[14'd4698] <= 32'h3e2bf262;
        mem[14'd4699] <= 32'h3e33ebf8;
        mem[14'd4700] <= 32'h3e480b9f;
        mem[14'd4701] <= 32'h3e3482be;
        mem[14'd4702] <= 32'hbd1a08d5;
        mem[14'd4703] <= 32'hbd5de418;
        mem[14'd4704] <= 32'hbcc36940;
        mem[14'd4705] <= 32'h3abd3427;
        mem[14'd4706] <= 32'h3c91164c;
        mem[14'd4707] <= 32'h3a1dc630;
        mem[14'd4708] <= 32'h3be4a013;
        mem[14'd4709] <= 32'hbc6aafca;
        mem[14'd4710] <= 32'hbabe2d21;
        mem[14'd4711] <= 32'h3b9264e8;
        mem[14'd4712] <= 32'hbca17f05;
        mem[14'd4713] <= 32'hbc8b4ade;
        mem[14'd4714] <= 32'hbcbe04d3;
        mem[14'd4715] <= 32'hbd69d7dc;
        mem[14'd4716] <= 32'hbdad3e01;
        mem[14'd4717] <= 32'hbb0b589d;
        mem[14'd4718] <= 32'hbc9d6344;
        mem[14'd4719] <= 32'h3d3a1d35;
        mem[14'd4720] <= 32'hbe02dbd7;
        mem[14'd4721] <= 32'hbe19884f;
        mem[14'd4722] <= 32'hbdb09aff;
        mem[14'd4723] <= 32'hbdd67af0;
        mem[14'd4724] <= 32'hbc27647b;
        mem[14'd4725] <= 32'hbdc905fa;
        mem[14'd4726] <= 32'hbcb19abe;
        mem[14'd4727] <= 32'h3d490bb9;
        mem[14'd4728] <= 32'h3d0426cc;
        mem[14'd4729] <= 32'h3d0a0038;
        mem[14'd4730] <= 32'hbb83cf87;
        mem[14'd4731] <= 32'hbc1e46c2;
        mem[14'd4732] <= 32'hbccadbe7;
        mem[14'd4733] <= 32'h3be7b89c;
        mem[14'd4734] <= 32'h3bc7fc05;
        mem[14'd4735] <= 32'h3cadc892;
        mem[14'd4736] <= 32'h3c2fd694;
        mem[14'd4737] <= 32'h3b264144;
        mem[14'd4738] <= 32'h3be6b854;
        mem[14'd4739] <= 32'h3c354039;
        mem[14'd4740] <= 32'hbc188438;
        mem[14'd4741] <= 32'hbcb4df6d;
        mem[14'd4742] <= 32'hbdc3e360;
        mem[14'd4743] <= 32'hbe2c692f;
        mem[14'd4744] <= 32'hbe6a5d95;
        mem[14'd4745] <= 32'hbe640e02;
        mem[14'd4746] <= 32'hbe3a9858;
        mem[14'd4747] <= 32'hbe877756;
        mem[14'd4748] <= 32'hbebf6857;
        mem[14'd4749] <= 32'hbe8dead5;
        mem[14'd4750] <= 32'hbe7cb5b7;
        mem[14'd4751] <= 32'hbe679f59;
        mem[14'd4752] <= 32'hbeadd5f8;
        mem[14'd4753] <= 32'hbec18e8b;
        mem[14'd4754] <= 32'hbe9a3098;
        mem[14'd4755] <= 32'hbe8d8bed;
        mem[14'd4756] <= 32'hbe17f469;
        mem[14'd4757] <= 32'hbdb9de5c;
        mem[14'd4758] <= 32'hbd5a780b;
        mem[14'd4759] <= 32'hbcf30808;
        mem[14'd4760] <= 32'hbc8da3a7;
        mem[14'd4761] <= 32'h3bb40177;
        mem[14'd4762] <= 32'hbc508c22;
        mem[14'd4763] <= 32'hbb960196;
        mem[14'd4764] <= 32'h3b92d7d8;
        mem[14'd4765] <= 32'hbc07e7db;
        mem[14'd4766] <= 32'h3c5ce497;
        mem[14'd4767] <= 32'h3c108b07;
        mem[14'd4768] <= 32'hbcc8933d;
        mem[14'd4769] <= 32'hbbac2642;
        mem[14'd4770] <= 32'hbd18dd95;
        mem[14'd4771] <= 32'hbd92b5b8;
        mem[14'd4772] <= 32'hbe0ec0b0;
        mem[14'd4773] <= 32'hbe473e73;
        mem[14'd4774] <= 32'hbe693081;
        mem[14'd4775] <= 32'hbe87fc32;
        mem[14'd4776] <= 32'hbe9139e6;
        mem[14'd4777] <= 32'hbea90307;
        mem[14'd4778] <= 32'hbecd0f43;
        mem[14'd4779] <= 32'hbeb2a078;
        mem[14'd4780] <= 32'hbe9a4eca;
        mem[14'd4781] <= 32'hbe94798b;
        mem[14'd4782] <= 32'hbe8c1262;
        mem[14'd4783] <= 32'hbe408771;
        mem[14'd4784] <= 32'hbdd064cc;
        mem[14'd4785] <= 32'hbd7337a1;
        mem[14'd4786] <= 32'hbca22f22;
        mem[14'd4787] <= 32'h3b224461;
        mem[14'd4788] <= 32'h3ac01775;
        mem[14'd4789] <= 32'h3c740b71;
        mem[14'd4790] <= 32'h3b5aec2b;
        mem[14'd4791] <= 32'h3c59c047;
        mem[14'd4792] <= 32'h3cbaeae5;
        mem[14'd4793] <= 32'hbaeae7a3;
        mem[14'd4794] <= 32'h3a91b684;
        mem[14'd4795] <= 32'hbb32261b;
        mem[14'd4796] <= 32'hbbf4ee7f;
        mem[14'd4797] <= 32'h3c60419e;
        mem[14'd4798] <= 32'h3b3ffc89;
        mem[14'd4799] <= 32'hbcaf9ff9;
        mem[14'd4800] <= 32'hbcc82b30;
        mem[14'd4801] <= 32'hbc1a1486;
        mem[14'd4802] <= 32'hbc84fa11;
        mem[14'd4803] <= 32'hbca8b893;
        mem[14'd4804] <= 32'hbcb82299;
        mem[14'd4805] <= 32'hbcd34ab9;
        mem[14'd4806] <= 32'hbd946d66;
        mem[14'd4807] <= 32'hbcd28826;
        mem[14'd4808] <= 32'hbc968aa4;
        mem[14'd4809] <= 32'hbd3c8955;
        mem[14'd4810] <= 32'hbd12fe50;
        mem[14'd4811] <= 32'hbcbd528c;
        mem[14'd4812] <= 32'hbca65010;
        mem[14'd4813] <= 32'hbcbb80d3;
        mem[14'd4814] <= 32'h3b843b27;
        mem[14'd4815] <= 32'hbca709bd;
        mem[14'd4816] <= 32'hbb5b3413;
        mem[14'd4817] <= 32'hbc041af9;
        mem[14'd4818] <= 32'hbc1e2a0e;
        mem[14'd4819] <= 32'h3bedda60;
        mem[14'd4820] <= 32'hbca52b8b;
        mem[14'd4821] <= 32'hbc7fadc5;
        mem[14'd4822] <= 32'h3c74a6d9;
        mem[14'd4823] <= 32'hbc0903c8;
        mem[14'd4824] <= 32'hbadc3d97;
        mem[14'd4825] <= 32'h3b9116bc;
        mem[14'd4826] <= 32'h3bbf3ad4;
        mem[14'd4827] <= 32'h39956381;
        mem[14'd4828] <= 32'hb9c40636;
        mem[14'd4829] <= 32'hbbdafc2a;
        mem[14'd4830] <= 32'h3c12ef79;
        mem[14'd4831] <= 32'hbbaa8064;
        mem[14'd4832] <= 32'h3bbc589b;
        mem[14'd4833] <= 32'h3abc3b79;
        mem[14'd4834] <= 32'h3aef812c;
        mem[14'd4835] <= 32'hbc030a46;
        mem[14'd4836] <= 32'h39e5cd03;
        mem[14'd4837] <= 32'h3b661fb5;
        mem[14'd4838] <= 32'hbb151ba0;
        mem[14'd4839] <= 32'hbb8b2f86;
        mem[14'd4840] <= 32'hbc186737;
        mem[14'd4841] <= 32'h3c24416d;
        mem[14'd4842] <= 32'h3ac2626e;
        mem[14'd4843] <= 32'h3c9052cd;
        mem[14'd4844] <= 32'h3a6592bb;
        mem[14'd4845] <= 32'h3bb3a6d2;
        mem[14'd4846] <= 32'hbc040539;
        mem[14'd4847] <= 32'hbb678299;
        mem[14'd4848] <= 32'h3b796c95;
        mem[14'd4849] <= 32'hbc0adcc8;
        mem[14'd4850] <= 32'hbbb3d415;
        mem[14'd4851] <= 32'h3a3a544c;
        mem[14'd4852] <= 32'h39809f38;
        mem[14'd4853] <= 32'h3b85132f;
        mem[14'd4854] <= 32'hbc7e1ded;
        mem[14'd4855] <= 32'h3b914f39;
        mem[14'd4856] <= 32'h3c20257c;
        mem[14'd4857] <= 32'h3b94b9f7;
        mem[14'd4858] <= 32'hbbc77dc4;
        mem[14'd4859] <= 32'h3b11cbb5;
        mem[14'd4860] <= 32'hbc842391;
        mem[14'd4861] <= 32'h3cca64ef;
        mem[14'd4862] <= 32'hbc08041b;
        mem[14'd4863] <= 32'h3a9debc8;
        mem[14'd4864] <= 32'h3b20df1b;
        mem[14'd4865] <= 32'hbaec94ee;
        mem[14'd4866] <= 32'h3c2dcb49;
        mem[14'd4867] <= 32'hbc2c22a6;
        mem[14'd4868] <= 32'h3c253bed;
        mem[14'd4869] <= 32'h3c3de56b;
        mem[14'd4870] <= 32'h3ad84440;
        mem[14'd4871] <= 32'hbba9808e;
        mem[14'd4872] <= 32'h3bc3982b;
        mem[14'd4873] <= 32'hbc41b5ea;
        mem[14'd4874] <= 32'h3c908fd7;
        mem[14'd4875] <= 32'hbc534666;
        mem[14'd4876] <= 32'h3c7ba052;
        mem[14'd4877] <= 32'hba963e26;
        mem[14'd4878] <= 32'hbbdd8c39;
        mem[14'd4879] <= 32'h3bbf40a7;
        mem[14'd4880] <= 32'hbb9d4cf0;
        mem[14'd4881] <= 32'hbc60b534;
        mem[14'd4882] <= 32'hbc62d79c;
        mem[14'd4883] <= 32'hbb2a32cf;
        mem[14'd4884] <= 32'hbc6d7d0b;
        mem[14'd4885] <= 32'hbbf54d1c;
        mem[14'd4886] <= 32'hbce66718;
        mem[14'd4887] <= 32'hbd49938a;
        mem[14'd4888] <= 32'hbd53c3ed;
        mem[14'd4889] <= 32'hbd80d386;
        mem[14'd4890] <= 32'hbd9dc75b;
        mem[14'd4891] <= 32'hbd4ec506;
        mem[14'd4892] <= 32'hbc5df3d6;
        mem[14'd4893] <= 32'h3ccb0079;
        mem[14'd4894] <= 32'h3c80077d;
        mem[14'd4895] <= 32'h3c635267;
        mem[14'd4896] <= 32'hbd19fa5c;
        mem[14'd4897] <= 32'hbcdc2900;
        mem[14'd4898] <= 32'hbcc1119d;
        mem[14'd4899] <= 32'hbc880080;
        mem[14'd4900] <= 32'h3b37958f;
        mem[14'd4901] <= 32'h3b3f1b44;
        mem[14'd4902] <= 32'h3b729a93;
        mem[14'd4903] <= 32'h3bb50bf9;
        mem[14'd4904] <= 32'h3c30f8b3;
        mem[14'd4905] <= 32'h3c0fd0e9;
        mem[14'd4906] <= 32'hbb91b71b;
        mem[14'd4907] <= 32'hbc758691;
        mem[14'd4908] <= 32'h3b52b123;
        mem[14'd4909] <= 32'hbc23d725;
        mem[14'd4910] <= 32'hbb5b5ce2;
        mem[14'd4911] <= 32'hbcc1c3c9;
        mem[14'd4912] <= 32'hbcf64e2d;
        mem[14'd4913] <= 32'hbd6de378;
        mem[14'd4914] <= 32'hbd36ffb7;
        mem[14'd4915] <= 32'hbdd35aa3;
        mem[14'd4916] <= 32'hbd6929d0;
        mem[14'd4917] <= 32'hbdb8c0af;
        mem[14'd4918] <= 32'hbd92e7a1;
        mem[14'd4919] <= 32'hbd09abf7;
        mem[14'd4920] <= 32'hbc458624;
        mem[14'd4921] <= 32'h3d8b9659;
        mem[14'd4922] <= 32'h3e0f74e5;
        mem[14'd4923] <= 32'h3e1619df;
        mem[14'd4924] <= 32'h3e215749;
        mem[14'd4925] <= 32'h3e0f484b;
        mem[14'd4926] <= 32'h3d9aa032;
        mem[14'd4927] <= 32'hbb2ed39d;
        mem[14'd4928] <= 32'h39929818;
        mem[14'd4929] <= 32'h3c8b07fe;
        mem[14'd4930] <= 32'h3c817d97;
        mem[14'd4931] <= 32'hbb8c9456;
        mem[14'd4932] <= 32'h3c8c9dfd;
        mem[14'd4933] <= 32'h3a8a3bb7;
        mem[14'd4934] <= 32'h3ca0246b;
        mem[14'd4935] <= 32'h3c60543a;
        mem[14'd4936] <= 32'hbd0fd73b;
        mem[14'd4937] <= 32'hbda98d81;
        mem[14'd4938] <= 32'hbdc744d1;
        mem[14'd4939] <= 32'hbe0b1f5a;
        mem[14'd4940] <= 32'hbe63ed03;
        mem[14'd4941] <= 32'hbe5672b8;
        mem[14'd4942] <= 32'hbdcd6e41;
        mem[14'd4943] <= 32'h3c14a4ef;
        mem[14'd4944] <= 32'hbd3469ae;
        mem[14'd4945] <= 32'hbe23f0d0;
        mem[14'd4946] <= 32'hbd05546a;
        mem[14'd4947] <= 32'h3e2f5184;
        mem[14'd4948] <= 32'h3df98dbc;
        mem[14'd4949] <= 32'h3e22d35a;
        mem[14'd4950] <= 32'h3e66ac75;
        mem[14'd4951] <= 32'h3dd23a87;
        mem[14'd4952] <= 32'hbd2b5ff6;
        mem[14'd4953] <= 32'h3e0b5500;
        mem[14'd4954] <= 32'h3ddbd6bc;
        mem[14'd4955] <= 32'h3e325d75;
        mem[14'd4956] <= 32'h3e3afa10;
        mem[14'd4957] <= 32'h3d7302ba;
        mem[14'd4958] <= 32'h3c7bc659;
        mem[14'd4959] <= 32'hbb7561a0;
        mem[14'd4960] <= 32'hbb25c069;
        mem[14'd4961] <= 32'h3c9e7651;
        mem[14'd4962] <= 32'h3a710d09;
        mem[14'd4963] <= 32'hbc594364;
        mem[14'd4964] <= 32'hbdb406f6;
        mem[14'd4965] <= 32'hbe1f6e00;
        mem[14'd4966] <= 32'hbe5e608e;
        mem[14'd4967] <= 32'hbe29b069;
        mem[14'd4968] <= 32'hbdd7c99e;
        mem[14'd4969] <= 32'h3c9e7f75;
        mem[14'd4970] <= 32'h3db2db86;
        mem[14'd4971] <= 32'h3d57cba5;
        mem[14'd4972] <= 32'hbd057be5;
        mem[14'd4973] <= 32'hbd5c6e61;
        mem[14'd4974] <= 32'hbde2a8fc;
        mem[14'd4975] <= 32'hbe0bfbd7;
        mem[14'd4976] <= 32'h3d212ce7;
        mem[14'd4977] <= 32'h3e135667;
        mem[14'd4978] <= 32'h3e0ef59a;
        mem[14'd4979] <= 32'h3cbfbbb7;
        mem[14'd4980] <= 32'h3e26a46a;
        mem[14'd4981] <= 32'h3dc28581;
        mem[14'd4982] <= 32'h3e7dc974;
        mem[14'd4983] <= 32'h3e842473;
        mem[14'd4984] <= 32'h3e8c8795;
        mem[14'd4985] <= 32'h3e27ad43;
        mem[14'd4986] <= 32'h3cecd914;
        mem[14'd4987] <= 32'hbc0aec94;
        mem[14'd4988] <= 32'h3b12576a;
        mem[14'd4989] <= 32'h3c2718d2;
        mem[14'd4990] <= 32'h3b80a005;
        mem[14'd4991] <= 32'hbda193a4;
        mem[14'd4992] <= 32'hbe301030;
        mem[14'd4993] <= 32'hbe2906d5;
        mem[14'd4994] <= 32'hbe0d7af8;
        mem[14'd4995] <= 32'hbcedf8cc;
        mem[14'd4996] <= 32'h3d743bee;
        mem[14'd4997] <= 32'h3cbb3ccf;
        mem[14'd4998] <= 32'h3c5c2e48;
        mem[14'd4999] <= 32'h3c82f1f3;
        mem[14'd5000] <= 32'h3ca0bfb4;
        mem[14'd5001] <= 32'hbd58ebfa;
        mem[14'd5002] <= 32'h3dc1ac47;
        mem[14'd5003] <= 32'hbd17b174;
        mem[14'd5004] <= 32'hbd85bd54;
        mem[14'd5005] <= 32'hbcb78b8f;
        mem[14'd5006] <= 32'h3d84024e;
        mem[14'd5007] <= 32'h3e35371e;
        mem[14'd5008] <= 32'h3e1679c1;
        mem[14'd5009] <= 32'h3bc419d4;
        mem[14'd5010] <= 32'h3e282a0e;
        mem[14'd5011] <= 32'h3ea971fd;
        mem[14'd5012] <= 32'h3f07f733;
        mem[14'd5013] <= 32'h3ea1abac;
        mem[14'd5014] <= 32'h3de7e44a;
        mem[14'd5015] <= 32'h3d07aa3e;
        mem[14'd5016] <= 32'h3c5f40d4;
        mem[14'd5017] <= 32'hbb20457d;
        mem[14'd5018] <= 32'h3b3839b7;
        mem[14'd5019] <= 32'hbdad37c8;
        mem[14'd5020] <= 32'hbe98b547;
        mem[14'd5021] <= 32'hbe5e2f77;
        mem[14'd5022] <= 32'hbdb37353;
        mem[14'd5023] <= 32'h3d0da157;
        mem[14'd5024] <= 32'h3e44ce16;
        mem[14'd5025] <= 32'h3dbb5b42;
        mem[14'd5026] <= 32'h3e2191ce;
        mem[14'd5027] <= 32'h3df9102e;
        mem[14'd5028] <= 32'h3d906314;
        mem[14'd5029] <= 32'hbdaa2848;
        mem[14'd5030] <= 32'h3dc7e615;
        mem[14'd5031] <= 32'hbdf03e5e;
        mem[14'd5032] <= 32'h3d8148fe;
        mem[14'd5033] <= 32'h3da1d643;
        mem[14'd5034] <= 32'h3d0f9d03;
        mem[14'd5035] <= 32'h3daffec1;
        mem[14'd5036] <= 32'h3ded92b6;
        mem[14'd5037] <= 32'h3de86084;
        mem[14'd5038] <= 32'h3e1dbd4c;
        mem[14'd5039] <= 32'h3eb86147;
        mem[14'd5040] <= 32'h3f236e6c;
        mem[14'd5041] <= 32'h3f08f631;
        mem[14'd5042] <= 32'h3e002d72;
        mem[14'd5043] <= 32'h3b699393;
        mem[14'd5044] <= 32'h3c86d601;
        mem[14'd5045] <= 32'hbc7daf6e;
        mem[14'd5046] <= 32'h3b07a8ae;
        mem[14'd5047] <= 32'hbdfe59b9;
        mem[14'd5048] <= 32'hbebb0cde;
        mem[14'd5049] <= 32'hbe82ce83;
        mem[14'd5050] <= 32'hbe0306c2;
        mem[14'd5051] <= 32'hbdc68581;
        mem[14'd5052] <= 32'h3df4a6c2;
        mem[14'd5053] <= 32'h3da2cfad;
        mem[14'd5054] <= 32'h3d95a08c;
        mem[14'd5055] <= 32'h3e190df2;
        mem[14'd5056] <= 32'h3c1e8a49;
        mem[14'd5057] <= 32'hbdc104da;
        mem[14'd5058] <= 32'hbe0397f2;
        mem[14'd5059] <= 32'hbe2faf8d;
        mem[14'd5060] <= 32'hbd75f930;
        mem[14'd5061] <= 32'hbc2c0527;
        mem[14'd5062] <= 32'hbcfaf76a;
        mem[14'd5063] <= 32'h3db1f265;
        mem[14'd5064] <= 32'h3e3ef579;
        mem[14'd5065] <= 32'h3e3108ba;
        mem[14'd5066] <= 32'h3e0d6fad;
        mem[14'd5067] <= 32'h3f08ce71;
        mem[14'd5068] <= 32'h3f603a00;
        mem[14'd5069] <= 32'h3f289dcc;
        mem[14'd5070] <= 32'h3e364af1;
        mem[14'd5071] <= 32'h3c99e218;
        mem[14'd5072] <= 32'hbb23527d;
        mem[14'd5073] <= 32'h3b837bbb;
        mem[14'd5074] <= 32'hbbd5e15b;
        mem[14'd5075] <= 32'hbde3ce51;
        mem[14'd5076] <= 32'hbe9029f3;
        mem[14'd5077] <= 32'hbe63a53a;
        mem[14'd5078] <= 32'hbd99a1d0;
        mem[14'd5079] <= 32'hbb4bdedf;
        mem[14'd5080] <= 32'h3e1a5fcc;
        mem[14'd5081] <= 32'h3d7fd137;
        mem[14'd5082] <= 32'h3e02e210;
        mem[14'd5083] <= 32'h3ea137cb;
        mem[14'd5084] <= 32'h3e1c3d08;
        mem[14'd5085] <= 32'hbd470194;
        mem[14'd5086] <= 32'hbe58d768;
        mem[14'd5087] <= 32'hbec0dbc3;
        mem[14'd5088] <= 32'hbeb8f379;
        mem[14'd5089] <= 32'hbe457777;
        mem[14'd5090] <= 32'hbd8502b4;
        mem[14'd5091] <= 32'hbda8f809;
        mem[14'd5092] <= 32'h3c8ebaef;
        mem[14'd5093] <= 32'h3e6fd866;
        mem[14'd5094] <= 32'h3e8556fb;
        mem[14'd5095] <= 32'h3f1110df;
        mem[14'd5096] <= 32'h3f8fbae2;
        mem[14'd5097] <= 32'h3f5604b0;
        mem[14'd5098] <= 32'h3e3bc137;
        mem[14'd5099] <= 32'h3c8b1061;
        mem[14'd5100] <= 32'h3be309b5;
        mem[14'd5101] <= 32'h3c6bcc3f;
        mem[14'd5102] <= 32'h391dfc5d;
        mem[14'd5103] <= 32'hbda796a7;
        mem[14'd5104] <= 32'hbe106698;
        mem[14'd5105] <= 32'hbe0273c6;
        mem[14'd5106] <= 32'hbc644efb;
        mem[14'd5107] <= 32'h3e225564;
        mem[14'd5108] <= 32'h3e898ecb;
        mem[14'd5109] <= 32'h3ea12a90;
        mem[14'd5110] <= 32'h3e8797c2;
        mem[14'd5111] <= 32'h3e86d912;
        mem[14'd5112] <= 32'h3e9a83b0;
        mem[14'd5113] <= 32'h3e5716d1;
        mem[14'd5114] <= 32'h3d526693;
        mem[14'd5115] <= 32'hbdf3c48e;
        mem[14'd5116] <= 32'hbe850ef0;
        mem[14'd5117] <= 32'hbebc5afd;
        mem[14'd5118] <= 32'hbeb18540;
        mem[14'd5119] <= 32'hbe9629f7;
        mem[14'd5120] <= 32'hbe2701d3;
        mem[14'd5121] <= 32'hbc893f1a;
        mem[14'd5122] <= 32'h3dc45866;
        mem[14'd5123] <= 32'h3f008c9f;
        mem[14'd5124] <= 32'h3f89767d;
        mem[14'd5125] <= 32'h3f6e70ce;
        mem[14'd5126] <= 32'h3e74b738;
        mem[14'd5127] <= 32'h3c779f18;
        mem[14'd5128] <= 32'h3b5c11a1;
        mem[14'd5129] <= 32'hbc7e2503;
        mem[14'd5130] <= 32'hbc225cfc;
        mem[14'd5131] <= 32'hbdb5adfb;
        mem[14'd5132] <= 32'hbd99fed7;
        mem[14'd5133] <= 32'hbc5af0ed;
        mem[14'd5134] <= 32'h3e42d331;
        mem[14'd5135] <= 32'h3dfba0c4;
        mem[14'd5136] <= 32'h3e36a56c;
        mem[14'd5137] <= 32'h3e08361d;
        mem[14'd5138] <= 32'h3e0ad451;
        mem[14'd5139] <= 32'h3e069925;
        mem[14'd5140] <= 32'h3e62cfe2;
        mem[14'd5141] <= 32'h3ecdd9a7;
        mem[14'd5142] <= 32'h3d9cc6f1;
        mem[14'd5143] <= 32'hbe1550d7;
        mem[14'd5144] <= 32'hbe28fe99;
        mem[14'd5145] <= 32'hbe573909;
        mem[14'd5146] <= 32'hbe53a084;
        mem[14'd5147] <= 32'hbeba7508;
        mem[14'd5148] <= 32'hbf10cd3a;
        mem[14'd5149] <= 32'hbeeb74ba;
        mem[14'd5150] <= 32'hbee5209f;
        mem[14'd5151] <= 32'hbd60b28d;
        mem[14'd5152] <= 32'h3eae8645;
        mem[14'd5153] <= 32'h3f01c8b5;
        mem[14'd5154] <= 32'h3e05f791;
        mem[14'd5155] <= 32'h3bba8cf6;
        mem[14'd5156] <= 32'hbc732755;
        mem[14'd5157] <= 32'h3b021f4a;
        mem[14'd5158] <= 32'hbc7a11a3;
        mem[14'd5159] <= 32'hbca6dcad;
        mem[14'd5160] <= 32'hbc6a8eaf;
        mem[14'd5161] <= 32'h3d184012;
        mem[14'd5162] <= 32'h3e6f5758;
        mem[14'd5163] <= 32'h3e002955;
        mem[14'd5164] <= 32'h3d0d73f7;
        mem[14'd5165] <= 32'hbccd8346;
        mem[14'd5166] <= 32'h3e5cc86b;
        mem[14'd5167] <= 32'h3e586c2c;
        mem[14'd5168] <= 32'h3e83e39c;
        mem[14'd5169] <= 32'h3e9c7fc6;
        mem[14'd5170] <= 32'hbd3a17c7;
        mem[14'd5171] <= 32'hbdd25c7f;
        mem[14'd5172] <= 32'hbea7a807;
        mem[14'd5173] <= 32'hbeb331d0;
        mem[14'd5174] <= 32'hbe8c1e16;
        mem[14'd5175] <= 32'hbea76c95;
        mem[14'd5176] <= 32'hbecf787b;
        mem[14'd5177] <= 32'hbf2f2511;
        mem[14'd5178] <= 32'hbf4ea877;
        mem[14'd5179] <= 32'hbf34b73d;
        mem[14'd5180] <= 32'hbefa1134;
        mem[14'd5181] <= 32'h3cc443c3;
        mem[14'd5182] <= 32'h3d42993b;
        mem[14'd5183] <= 32'hbccce28d;
        mem[14'd5184] <= 32'hbb5ef0e9;
        mem[14'd5185] <= 32'h3adee320;
        mem[14'd5186] <= 32'h3bb674df;
        mem[14'd5187] <= 32'hbbc9f0de;
        mem[14'd5188] <= 32'h3d3f07e2;
        mem[14'd5189] <= 32'h3da01e64;
        mem[14'd5190] <= 32'h3d136d0b;
        mem[14'd5191] <= 32'h3e17613a;
        mem[14'd5192] <= 32'h3d0a5fa0;
        mem[14'd5193] <= 32'h3d8b9695;
        mem[14'd5194] <= 32'h3e5bbff1;
        mem[14'd5195] <= 32'h3e9cddca;
        mem[14'd5196] <= 32'h3eb27142;
        mem[14'd5197] <= 32'h3e5aa526;
        mem[14'd5198] <= 32'hbce1a80d;
        mem[14'd5199] <= 32'hbe7e4866;
        mem[14'd5200] <= 32'hbee9aef1;
        mem[14'd5201] <= 32'hbe708baa;
        mem[14'd5202] <= 32'hbe125ad8;
        mem[14'd5203] <= 32'hbd91c784;
        mem[14'd5204] <= 32'hbdbb4d8e;
        mem[14'd5205] <= 32'hbe90e9d0;
        mem[14'd5206] <= 32'hbec67f4d;
        mem[14'd5207] <= 32'hbf0bb202;
        mem[14'd5208] <= 32'hbee0dfcc;
        mem[14'd5209] <= 32'hbdb1350b;
        mem[14'd5210] <= 32'h3a87e483;
        mem[14'd5211] <= 32'h3c430f2e;
        mem[14'd5212] <= 32'h3c0b3a4b;
        mem[14'd5213] <= 32'hbbb4ac99;
        mem[14'd5214] <= 32'hbc0f7bc1;
        mem[14'd5215] <= 32'h3c74746c;
        mem[14'd5216] <= 32'h3d1490c5;
        mem[14'd5217] <= 32'hbd363417;
        mem[14'd5218] <= 32'hbd2a3c38;
        mem[14'd5219] <= 32'h3a0df4fe;
        mem[14'd5220] <= 32'h3d6a1b7a;
        mem[14'd5221] <= 32'h3e28fc50;
        mem[14'd5222] <= 32'h3e8e99aa;
        mem[14'd5223] <= 32'h3d07ccf1;
        mem[14'd5224] <= 32'h3db6ef6a;
        mem[14'd5225] <= 32'h3d01533f;
        mem[14'd5226] <= 32'hbd91031d;
        mem[14'd5227] <= 32'hbe36a870;
        mem[14'd5228] <= 32'hbe83db79;
        mem[14'd5229] <= 32'hbe75db17;
        mem[14'd5230] <= 32'hbe2c0f71;
        mem[14'd5231] <= 32'hbe574b4d;
        mem[14'd5232] <= 32'hbda33294;
        mem[14'd5233] <= 32'hbe067cdb;
        mem[14'd5234] <= 32'hbd449f9e;
        mem[14'd5235] <= 32'hbe47a159;
        mem[14'd5236] <= 32'hbe30f60d;
        mem[14'd5237] <= 32'hbdd8c4a7;
        mem[14'd5238] <= 32'hbcb4875c;
        mem[14'd5239] <= 32'h3c10821f;
        mem[14'd5240] <= 32'h3a9159dd;
        mem[14'd5241] <= 32'h3a5f0597;
        mem[14'd5242] <= 32'hbc4e991e;
        mem[14'd5243] <= 32'h3b8b8ef2;
        mem[14'd5244] <= 32'hbd23613f;
        mem[14'd5245] <= 32'hbe382605;
        mem[14'd5246] <= 32'hbe0b736a;
        mem[14'd5247] <= 32'hbe497d45;
        mem[14'd5248] <= 32'hbb0e59c7;
        mem[14'd5249] <= 32'h3e0a0cc4;
        mem[14'd5250] <= 32'h3e21986d;
        mem[14'd5251] <= 32'h3d7f5589;
        mem[14'd5252] <= 32'h3dec5341;
        mem[14'd5253] <= 32'hbd5be867;
        mem[14'd5254] <= 32'hbe8568a8;
        mem[14'd5255] <= 32'hbe84b9f4;
        mem[14'd5256] <= 32'hbe3e2058;
        mem[14'd5257] <= 32'hbe644e7d;
        mem[14'd5258] <= 32'h3dce4d27;
        mem[14'd5259] <= 32'hbd76449b;
        mem[14'd5260] <= 32'hbde8005d;
        mem[14'd5261] <= 32'hbcd0d526;
        mem[14'd5262] <= 32'hbd84896e;
        mem[14'd5263] <= 32'h3a8f9d31;
        mem[14'd5264] <= 32'hbce89fa5;
        mem[14'd5265] <= 32'hbd7baa0d;
        mem[14'd5266] <= 32'hbd13a905;
        mem[14'd5267] <= 32'hbbf01972;
        mem[14'd5268] <= 32'hbc5facc1;
        mem[14'd5269] <= 32'hba5407e1;
        mem[14'd5270] <= 32'hbb00ca1d;
        mem[14'd5271] <= 32'hbc8ec329;
        mem[14'd5272] <= 32'hbd776f26;
        mem[14'd5273] <= 32'hbe1f19b8;
        mem[14'd5274] <= 32'hbe3772e8;
        mem[14'd5275] <= 32'hbebd8d18;
        mem[14'd5276] <= 32'hbe964ba9;
        mem[14'd5277] <= 32'hbe8cfe32;
        mem[14'd5278] <= 32'hbdfc6bab;
        mem[14'd5279] <= 32'hbe04ca7c;
        mem[14'd5280] <= 32'hbd05f110;
        mem[14'd5281] <= 32'hbda068e8;
        mem[14'd5282] <= 32'hbe87e5b0;
        mem[14'd5283] <= 32'hbe19c277;
        mem[14'd5284] <= 32'hbe768bb1;
        mem[14'd5285] <= 32'hbdf10cb0;
        mem[14'd5286] <= 32'hbdcf56df;
        mem[14'd5287] <= 32'hbc7f2aa8;
        mem[14'd5288] <= 32'h3d0850c7;
        mem[14'd5289] <= 32'hba57f032;
        mem[14'd5290] <= 32'h3dbe6b17;
        mem[14'd5291] <= 32'h3dae0c1d;
        mem[14'd5292] <= 32'h3c85ed4f;
        mem[14'd5293] <= 32'hbd837bc7;
        mem[14'd5294] <= 32'hbd0eb247;
        mem[14'd5295] <= 32'hbc0e7d0e;
        mem[14'd5296] <= 32'hbb182db4;
        mem[14'd5297] <= 32'h3ccbef28;
        mem[14'd5298] <= 32'hbc5cdcc4;
        mem[14'd5299] <= 32'h3c920423;
        mem[14'd5300] <= 32'h3cb1e567;
        mem[14'd5301] <= 32'h3de22cfd;
        mem[14'd5302] <= 32'h3e80c266;
        mem[14'd5303] <= 32'hbe4cbb6a;
        mem[14'd5304] <= 32'hbe982d6a;
        mem[14'd5305] <= 32'hbe9bcb6b;
        mem[14'd5306] <= 32'hbe9a7b2a;
        mem[14'd5307] <= 32'hbe87f062;
        mem[14'd5308] <= 32'hbed31aa1;
        mem[14'd5309] <= 32'hbed06697;
        mem[14'd5310] <= 32'hbea112af;
        mem[14'd5311] <= 32'hbda989bf;
        mem[14'd5312] <= 32'h3cdf75ef;
        mem[14'd5313] <= 32'h3dc16637;
        mem[14'd5314] <= 32'h3e247ec0;
        mem[14'd5315] <= 32'h3cc47347;
        mem[14'd5316] <= 32'h3dbbd734;
        mem[14'd5317] <= 32'h3da013ae;
        mem[14'd5318] <= 32'h3bf5b02a;
        mem[14'd5319] <= 32'h3de4d9e9;
        mem[14'd5320] <= 32'h3d84d841;
        mem[14'd5321] <= 32'hbd81d712;
        mem[14'd5322] <= 32'hbc5826be;
        mem[14'd5323] <= 32'hbc5e8a0f;
        mem[14'd5324] <= 32'hbc50fe3a;
        mem[14'd5325] <= 32'h3c4c3c9d;
        mem[14'd5326] <= 32'hbd1d8200;
        mem[14'd5327] <= 32'h3c69a2b2;
        mem[14'd5328] <= 32'h3e28b237;
        mem[14'd5329] <= 32'h3e81d916;
        mem[14'd5330] <= 32'h3ee7688d;
        mem[14'd5331] <= 32'h3e463258;
        mem[14'd5332] <= 32'hbd0f6774;
        mem[14'd5333] <= 32'hbe09a1ee;
        mem[14'd5334] <= 32'hbe2f8b42;
        mem[14'd5335] <= 32'hbdfb28df;
        mem[14'd5336] <= 32'hbe35704c;
        mem[14'd5337] <= 32'hbd928c61;
        mem[14'd5338] <= 32'hbc0742bf;
        mem[14'd5339] <= 32'hbc2479b1;
        mem[14'd5340] <= 32'h3c1d172f;
        mem[14'd5341] <= 32'h3e0921a3;
        mem[14'd5342] <= 32'hbc6fb78c;
        mem[14'd5343] <= 32'h3d69ba43;
        mem[14'd5344] <= 32'h3db53c76;
        mem[14'd5345] <= 32'h3d61efd2;
        mem[14'd5346] <= 32'h3d906df4;
        mem[14'd5347] <= 32'h3dff16b0;
        mem[14'd5348] <= 32'h3e097c03;
        mem[14'd5349] <= 32'hbd047471;
        mem[14'd5350] <= 32'hbc83ba87;
        mem[14'd5351] <= 32'hbc22a67e;
        mem[14'd5352] <= 32'h3c153b75;
        mem[14'd5353] <= 32'h3c386fd6;
        mem[14'd5354] <= 32'h3c17ea7e;
        mem[14'd5355] <= 32'h3d29310a;
        mem[14'd5356] <= 32'h3e6008f5;
        mem[14'd5357] <= 32'h3e4d1e4d;
        mem[14'd5358] <= 32'h3eb6dd92;
        mem[14'd5359] <= 32'h3e3c2825;
        mem[14'd5360] <= 32'h3e903a81;
        mem[14'd5361] <= 32'h3dc72cf5;
        mem[14'd5362] <= 32'h3cee8d27;
        mem[14'd5363] <= 32'h3da8467e;
        mem[14'd5364] <= 32'h3d29d789;
        mem[14'd5365] <= 32'h3d9c818e;
        mem[14'd5366] <= 32'h3c64f454;
        mem[14'd5367] <= 32'h3cb85538;
        mem[14'd5368] <= 32'hbd7eb232;
        mem[14'd5369] <= 32'hbd4e7b13;
        mem[14'd5370] <= 32'h3d59aa6c;
        mem[14'd5371] <= 32'h3d2a7b5b;
        mem[14'd5372] <= 32'h3e0d8bb7;
        mem[14'd5373] <= 32'h3dc5a869;
        mem[14'd5374] <= 32'h3e10bdf6;
        mem[14'd5375] <= 32'h3e379b19;
        mem[14'd5376] <= 32'h3e1562e0;
        mem[14'd5377] <= 32'hbc5265f9;
        mem[14'd5378] <= 32'hbc947915;
        mem[14'd5379] <= 32'h3b5e8234;
        mem[14'd5380] <= 32'hbb6a278e;
        mem[14'd5381] <= 32'hba1786d9;
        mem[14'd5382] <= 32'h3b762fb6;
        mem[14'd5383] <= 32'h3d505906;
        mem[14'd5384] <= 32'h3dfa597b;
        mem[14'd5385] <= 32'h3e819317;
        mem[14'd5386] <= 32'h3e29f908;
        mem[14'd5387] <= 32'h3c0ae778;
        mem[14'd5388] <= 32'h3e769a80;
        mem[14'd5389] <= 32'h3e5b51c6;
        mem[14'd5390] <= 32'h3d38094f;
        mem[14'd5391] <= 32'h3e0346ec;
        mem[14'd5392] <= 32'h3d06d42c;
        mem[14'd5393] <= 32'h3d6c173c;
        mem[14'd5394] <= 32'hbd431073;
        mem[14'd5395] <= 32'hbc7a9741;
        mem[14'd5396] <= 32'h3dd1dc16;
        mem[14'd5397] <= 32'h3e12153d;
        mem[14'd5398] <= 32'h3da03b42;
        mem[14'd5399] <= 32'h3d9e2fe5;
        mem[14'd5400] <= 32'h3c3141e9;
        mem[14'd5401] <= 32'h3da78729;
        mem[14'd5402] <= 32'h3e9cb680;
        mem[14'd5403] <= 32'h3e4731a0;
        mem[14'd5404] <= 32'h3d9a8e0e;
        mem[14'd5405] <= 32'h3cb0c19b;
        mem[14'd5406] <= 32'hbbdb47e4;
        mem[14'd5407] <= 32'h3c33d6e6;
        mem[14'd5408] <= 32'hbbb4d856;
        mem[14'd5409] <= 32'h3c745f37;
        mem[14'd5410] <= 32'hbc1f50df;
        mem[14'd5411] <= 32'h3aaca014;
        mem[14'd5412] <= 32'h3e17e2b9;
        mem[14'd5413] <= 32'h3de6553c;
        mem[14'd5414] <= 32'h3ded8fb9;
        mem[14'd5415] <= 32'h3e192fe8;
        mem[14'd5416] <= 32'h3e36f4e1;
        mem[14'd5417] <= 32'h3df85096;
        mem[14'd5418] <= 32'h3d7de45b;
        mem[14'd5419] <= 32'h3e1562a3;
        mem[14'd5420] <= 32'h3dd057d7;
        mem[14'd5421] <= 32'h3d8975c4;
        mem[14'd5422] <= 32'h3ddf9bd0;
        mem[14'd5423] <= 32'h3dc2e89e;
        mem[14'd5424] <= 32'h3ce3a78b;
        mem[14'd5425] <= 32'h3d8b0e17;
        mem[14'd5426] <= 32'hbc5fc65a;
        mem[14'd5427] <= 32'h3c9bfee8;
        mem[14'd5428] <= 32'h3e1d6338;
        mem[14'd5429] <= 32'h3e94ecda;
        mem[14'd5430] <= 32'h3e9d2395;
        mem[14'd5431] <= 32'h3e3d83a6;
        mem[14'd5432] <= 32'h3d9ffdc0;
        mem[14'd5433] <= 32'h3ce714b0;
        mem[14'd5434] <= 32'h3c03e739;
        mem[14'd5435] <= 32'hbc86079d;
        mem[14'd5436] <= 32'h3a8a98f5;
        mem[14'd5437] <= 32'hbbf1b86e;
        mem[14'd5438] <= 32'hba8332f6;
        mem[14'd5439] <= 32'hbb62889b;
        mem[14'd5440] <= 32'h3e08a6a4;
        mem[14'd5441] <= 32'hbd196c3b;
        mem[14'd5442] <= 32'hbe0010f5;
        mem[14'd5443] <= 32'hbc1dfb72;
        mem[14'd5444] <= 32'h3cf95c1c;
        mem[14'd5445] <= 32'h3d4564fc;
        mem[14'd5446] <= 32'hbd7a6d6c;
        mem[14'd5447] <= 32'h3d88007e;
        mem[14'd5448] <= 32'h3e2f7b9e;
        mem[14'd5449] <= 32'h3e59387b;
        mem[14'd5450] <= 32'h3e0444c3;
        mem[14'd5451] <= 32'h3d6a9b13;
        mem[14'd5452] <= 32'h3e029f93;
        mem[14'd5453] <= 32'h3d40d16b;
        mem[14'd5454] <= 32'h3dd9c986;
        mem[14'd5455] <= 32'h3de19d19;
        mem[14'd5456] <= 32'h3e0bf54c;
        mem[14'd5457] <= 32'h3df85582;
        mem[14'd5458] <= 32'h3e281659;
        mem[14'd5459] <= 32'h3e12ccd6;
        mem[14'd5460] <= 32'h3d87b27d;
        mem[14'd5461] <= 32'h3d0f6024;
        mem[14'd5462] <= 32'h3cc3e9e7;
        mem[14'd5463] <= 32'hbc73ef1f;
        mem[14'd5464] <= 32'h3a68980b;
        mem[14'd5465] <= 32'hbbae10fd;
        mem[14'd5466] <= 32'hbbc7d877;
        mem[14'd5467] <= 32'h3c7f0126;
        mem[14'd5468] <= 32'h3d838fce;
        mem[14'd5469] <= 32'h3db9be4c;
        mem[14'd5470] <= 32'hbd10a192;
        mem[14'd5471] <= 32'hbe031f57;
        mem[14'd5472] <= 32'h3dc7a7bb;
        mem[14'd5473] <= 32'h3de9cd28;
        mem[14'd5474] <= 32'h3e427afa;
        mem[14'd5475] <= 32'h3dd92a2c;
        mem[14'd5476] <= 32'h3df9c661;
        mem[14'd5477] <= 32'hbcd90cc1;
        mem[14'd5478] <= 32'h3db046e0;
        mem[14'd5479] <= 32'h3d20bb63;
        mem[14'd5480] <= 32'h3e03b559;
        mem[14'd5481] <= 32'hbc4b5b44;
        mem[14'd5482] <= 32'hbe0f54a1;
        mem[14'd5483] <= 32'hbc4be114;
        mem[14'd5484] <= 32'h3d4cbe74;
        mem[14'd5485] <= 32'h3cfd6ad1;
        mem[14'd5486] <= 32'h3d8a3954;
        mem[14'd5487] <= 32'h3d980022;
        mem[14'd5488] <= 32'h3d706a70;
        mem[14'd5489] <= 32'hbb920921;
        mem[14'd5490] <= 32'hba3fdb95;
        mem[14'd5491] <= 32'hb994e463;
        mem[14'd5492] <= 32'h3c0a57d5;
        mem[14'd5493] <= 32'hbcc5de75;
        mem[14'd5494] <= 32'h3a2cb695;
        mem[14'd5495] <= 32'h3c269dc3;
        mem[14'd5496] <= 32'hbc823bd3;
        mem[14'd5497] <= 32'hbba5a39a;
        mem[14'd5498] <= 32'hbcacf80f;
        mem[14'd5499] <= 32'h3bddc877;
        mem[14'd5500] <= 32'h3d91d9d4;
        mem[14'd5501] <= 32'h3e8babe8;
        mem[14'd5502] <= 32'h3e4731fb;
        mem[14'd5503] <= 32'h3e355210;
        mem[14'd5504] <= 32'h3e644b6a;
        mem[14'd5505] <= 32'h3e8b94f2;
        mem[14'd5506] <= 32'h3e884cea;
        mem[14'd5507] <= 32'h3e599997;
        mem[14'd5508] <= 32'h3dd31814;
        mem[14'd5509] <= 32'h3e21ce24;
        mem[14'd5510] <= 32'h3de78064;
        mem[14'd5511] <= 32'h3d0fdb7e;
        mem[14'd5512] <= 32'h3d218a16;
        mem[14'd5513] <= 32'h3c3a85ef;
        mem[14'd5514] <= 32'h3d90a867;
        mem[14'd5515] <= 32'h3d5cacbe;
        mem[14'd5516] <= 32'h3ce58480;
        mem[14'd5517] <= 32'h3b19f7d0;
        mem[14'd5518] <= 32'h3abc2ba6;
        mem[14'd5519] <= 32'hbb4ba914;
        mem[14'd5520] <= 32'hbc5d5817;
        mem[14'd5521] <= 32'hbbc45d62;
        mem[14'd5522] <= 32'hbb7f5a43;
        mem[14'd5523] <= 32'h3c2b431b;
        mem[14'd5524] <= 32'h3c930ac4;
        mem[14'd5525] <= 32'hbbf5ce9e;
        mem[14'd5526] <= 32'hbc9a3cb0;
        mem[14'd5527] <= 32'hbd07602b;
        mem[14'd5528] <= 32'h3bc1033a;
        mem[14'd5529] <= 32'h3ddd2ab3;
        mem[14'd5530] <= 32'h3e02433f;
        mem[14'd5531] <= 32'h3e37c6f2;
        mem[14'd5532] <= 32'h3e502ec9;
        mem[14'd5533] <= 32'h3e5753e8;
        mem[14'd5534] <= 32'h3df17ed5;
        mem[14'd5535] <= 32'h3e6f00a7;
        mem[14'd5536] <= 32'h3e42cdd6;
        mem[14'd5537] <= 32'h3e338fe0;
        mem[14'd5538] <= 32'h3dab5e0e;
        mem[14'd5539] <= 32'h3d6eeac3;
        mem[14'd5540] <= 32'h3cac4205;
        mem[14'd5541] <= 32'h3d574c75;
        mem[14'd5542] <= 32'h3dc26e97;
        mem[14'd5543] <= 32'h3d8ab9f9;
        mem[14'd5544] <= 32'h3d288bb3;
        mem[14'd5545] <= 32'h3cc3b1c0;
        mem[14'd5546] <= 32'h3c6168f6;
        mem[14'd5547] <= 32'h3c178899;
        mem[14'd5548] <= 32'hbbf8af0a;
        mem[14'd5549] <= 32'h38707f9b;
        mem[14'd5550] <= 32'h3c6e81a0;
        mem[14'd5551] <= 32'hbc250053;
        mem[14'd5552] <= 32'hbc071140;
        mem[14'd5553] <= 32'hbb609544;
        mem[14'd5554] <= 32'h3b4ac96e;
        mem[14'd5555] <= 32'hbd321f9e;
        mem[14'd5556] <= 32'hbd9d5ec4;
        mem[14'd5557] <= 32'hbd00eee6;
        mem[14'd5558] <= 32'h3a2cdbe0;
        mem[14'd5559] <= 32'h3d11aff1;
        mem[14'd5560] <= 32'h3d11452b;
        mem[14'd5561] <= 32'h3c0ba28c;
        mem[14'd5562] <= 32'hbd054082;
        mem[14'd5563] <= 32'h3ccb73d4;
        mem[14'd5564] <= 32'h3b581602;
        mem[14'd5565] <= 32'hbd2698e2;
        mem[14'd5566] <= 32'hbd63680c;
        mem[14'd5567] <= 32'hbc6e7de6;
        mem[14'd5568] <= 32'hbbebfd29;
        mem[14'd5569] <= 32'h3c322384;
        mem[14'd5570] <= 32'h3c98b9fb;
        mem[14'd5571] <= 32'h3bc2a5aa;
        mem[14'd5572] <= 32'h3c87973e;
        mem[14'd5573] <= 32'hbc0b4d61;
        mem[14'd5574] <= 32'h3c737f4c;
        mem[14'd5575] <= 32'hbc2ce052;
        mem[14'd5576] <= 32'hbaf2f28f;
        mem[14'd5577] <= 32'hbbab86e0;
        mem[14'd5578] <= 32'h3b9a3767;
        mem[14'd5579] <= 32'hbc1c6730;
        mem[14'd5580] <= 32'hbb8111a3;
        mem[14'd5581] <= 32'h3b9d56e4;
        mem[14'd5582] <= 32'hbb00a58e;
        mem[14'd5583] <= 32'h3c234416;
        mem[14'd5584] <= 32'hba86500b;
        mem[14'd5585] <= 32'h3bef91a4;
        mem[14'd5586] <= 32'h3c9c5611;
        mem[14'd5587] <= 32'hbc265dea;
        mem[14'd5588] <= 32'h3c0a830d;
        mem[14'd5589] <= 32'hbb6bbd3c;
        mem[14'd5590] <= 32'hbc3bab58;
        mem[14'd5591] <= 32'hbc7019e7;
        mem[14'd5592] <= 32'hbc8ec5a3;
        mem[14'd5593] <= 32'hbcaa8133;
        mem[14'd5594] <= 32'hbc9052eb;
        mem[14'd5595] <= 32'hbc21fbb2;
        mem[14'd5596] <= 32'hbb8ccbaf;
        mem[14'd5597] <= 32'hbc8dcda5;
        mem[14'd5598] <= 32'hbc10d380;
        mem[14'd5599] <= 32'hbb1aa63a;
        mem[14'd5600] <= 32'h3c213b84;
        mem[14'd5601] <= 32'h3b9f61e0;
        mem[14'd5602] <= 32'h3c2c3993;
        mem[14'd5603] <= 32'h3b775ade;
        mem[14'd5604] <= 32'hbbab9653;
        mem[14'd5605] <= 32'h3b1ca4b8;
        mem[14'd5606] <= 32'h3be3de20;
        mem[14'd5607] <= 32'hbaff5dbc;
        mem[14'd5608] <= 32'hbc69f9b5;
        mem[14'd5609] <= 32'hbacc61cd;
        mem[14'd5610] <= 32'h3beaef93;
        mem[14'd5611] <= 32'hb92bf2cc;
        mem[14'd5612] <= 32'hb9149615;
        mem[14'd5613] <= 32'hbb44c98f;
        mem[14'd5614] <= 32'hbbceffe2;
        mem[14'd5615] <= 32'hbb1bc2d3;
        mem[14'd5616] <= 32'hba871266;
        mem[14'd5617] <= 32'hbbc3758e;
        mem[14'd5618] <= 32'h3c372a44;
        mem[14'd5619] <= 32'h39f44776;
        mem[14'd5620] <= 32'h3b85ce07;
        mem[14'd5621] <= 32'hbba6c650;
        mem[14'd5622] <= 32'h3c2fad3e;
        mem[14'd5623] <= 32'h3c3d5559;
        mem[14'd5624] <= 32'h3b376dfe;
        mem[14'd5625] <= 32'hbb8ed35c;
        mem[14'd5626] <= 32'h3c515793;
        mem[14'd5627] <= 32'h3bef6134;
        mem[14'd5628] <= 32'hbb1f2f67;
        mem[14'd5629] <= 32'h3b965ca2;
        mem[14'd5630] <= 32'hba41e359;
        mem[14'd5631] <= 32'hbc2f48c6;
        mem[14'd5632] <= 32'h3bd0c342;
        mem[14'd5633] <= 32'hba552477;
        mem[14'd5634] <= 32'hbc8f6b81;
        mem[14'd5635] <= 32'hbbe68d32;
        mem[14'd5636] <= 32'hbb5f595f;
        mem[14'd5637] <= 32'h3c0bc991;
        mem[14'd5638] <= 32'h3cc0eb23;
        mem[14'd5639] <= 32'h3d20c121;
        mem[14'd5640] <= 32'h3cfa5c63;
        mem[14'd5641] <= 32'h3d3f67b6;
        mem[14'd5642] <= 32'h3d26892a;
        mem[14'd5643] <= 32'h3d8ffe76;
        mem[14'd5644] <= 32'h3db0ccec;
        mem[14'd5645] <= 32'h3d73286e;
        mem[14'd5646] <= 32'h3d04d817;
        mem[14'd5647] <= 32'h3d000c9c;
        mem[14'd5648] <= 32'h3c413fcf;
        mem[14'd5649] <= 32'h3c716ecb;
        mem[14'd5650] <= 32'h3c9126c7;
        mem[14'd5651] <= 32'h3d1dc3d0;
        mem[14'd5652] <= 32'h3bab447c;
        mem[14'd5653] <= 32'h3c5afadd;
        mem[14'd5654] <= 32'h3c9a614a;
        mem[14'd5655] <= 32'hbc234321;
        mem[14'd5656] <= 32'hbbfe85f9;
        mem[14'd5657] <= 32'h3ca450b0;
        mem[14'd5658] <= 32'hbce245c7;
        mem[14'd5659] <= 32'hb9b0c989;
        mem[14'd5660] <= 32'h3b1398ef;
        mem[14'd5661] <= 32'h3bc0e367;
        mem[14'd5662] <= 32'hba806d7d;
        mem[14'd5663] <= 32'hbbb83837;
        mem[14'd5664] <= 32'h3bcc8b59;
        mem[14'd5665] <= 32'h3b99ec43;
        mem[14'd5666] <= 32'h3d26efd1;
        mem[14'd5667] <= 32'h3d8dd6e1;
        mem[14'd5668] <= 32'h3dedabb4;
        mem[14'd5669] <= 32'h3dd98524;
        mem[14'd5670] <= 32'h3e62f0b6;
        mem[14'd5671] <= 32'h3e79edaf;
        mem[14'd5672] <= 32'h3e8b711d;
        mem[14'd5673] <= 32'h3e87ac19;
        mem[14'd5674] <= 32'h3e60f6f0;
        mem[14'd5675] <= 32'h3e40d167;
        mem[14'd5676] <= 32'h3e2e2172;
        mem[14'd5677] <= 32'h3e3a2085;
        mem[14'd5678] <= 32'h3e315ae6;
        mem[14'd5679] <= 32'h3e33c299;
        mem[14'd5680] <= 32'h3dfff5fe;
        mem[14'd5681] <= 32'h3dd3b2df;
        mem[14'd5682] <= 32'h3dc9d350;
        mem[14'd5683] <= 32'h3d3cd4e2;
        mem[14'd5684] <= 32'hbb60bab4;
        mem[14'd5685] <= 32'hbb7e05a1;
        mem[14'd5686] <= 32'hbc207234;
        mem[14'd5687] <= 32'h3b6eeeeb;
        mem[14'd5688] <= 32'hbc4d0907;
        mem[14'd5689] <= 32'h3ba7b6a6;
        mem[14'd5690] <= 32'h3bcec270;
        mem[14'd5691] <= 32'h3c158841;
        mem[14'd5692] <= 32'h3c6e2857;
        mem[14'd5693] <= 32'h3bab01a6;
        mem[14'd5694] <= 32'h3d7a6d58;
        mem[14'd5695] <= 32'h3da8acac;
        mem[14'd5696] <= 32'h3e00120e;
        mem[14'd5697] <= 32'h3e16a5e5;
        mem[14'd5698] <= 32'h3e4a371b;
        mem[14'd5699] <= 32'h3e7f37a2;
        mem[14'd5700] <= 32'h3e37d73c;
        mem[14'd5701] <= 32'h3e6ef9af;
        mem[14'd5702] <= 32'h3e445a31;
        mem[14'd5703] <= 32'h3e259b87;
        mem[14'd5704] <= 32'h3dc97b60;
        mem[14'd5705] <= 32'h3dc2a5cf;
        mem[14'd5706] <= 32'h3e432e22;
        mem[14'd5707] <= 32'h3e6da9ef;
        mem[14'd5708] <= 32'h3dfcfba7;
        mem[14'd5709] <= 32'h3e1dd391;
        mem[14'd5710] <= 32'h3e274de0;
        mem[14'd5711] <= 32'h3e12874a;
        mem[14'd5712] <= 32'h3d966e7b;
        mem[14'd5713] <= 32'hbbea42d1;
        mem[14'd5714] <= 32'h3ba6806a;
        mem[14'd5715] <= 32'h3afd4f38;
        mem[14'd5716] <= 32'hbcabf9f6;
        mem[14'd5717] <= 32'hbc245b1a;
        mem[14'd5718] <= 32'hbc1ec379;
        mem[14'd5719] <= 32'hb9aaec8d;
        mem[14'd5720] <= 32'hbc857928;
        mem[14'd5721] <= 32'h3b50df43;
        mem[14'd5722] <= 32'h3bcef443;
        mem[14'd5723] <= 32'h3d12827b;
        mem[14'd5724] <= 32'h3da02f4a;
        mem[14'd5725] <= 32'h3cc6c50f;
        mem[14'd5726] <= 32'h3d879b80;
        mem[14'd5727] <= 32'hbd22230e;
        mem[14'd5728] <= 32'hbdebac24;
        mem[14'd5729] <= 32'hbd8367a9;
        mem[14'd5730] <= 32'hbd9b4e3a;
        mem[14'd5731] <= 32'hbdf49b44;
        mem[14'd5732] <= 32'h3d2fdee9;
        mem[14'd5733] <= 32'h3dc2d8c6;
        mem[14'd5734] <= 32'h3d528f4f;
        mem[14'd5735] <= 32'h3ded930d;
        mem[14'd5736] <= 32'h3e58343c;
        mem[14'd5737] <= 32'h3e63e388;
        mem[14'd5738] <= 32'h3e8a8dab;
        mem[14'd5739] <= 32'h3e39040c;
        mem[14'd5740] <= 32'h3b9864fc;
        mem[14'd5741] <= 32'hbc83c6ae;
        mem[14'd5742] <= 32'h3aeed399;
        mem[14'd5743] <= 32'h3c44a327;
        mem[14'd5744] <= 32'hba14ec68;
        mem[14'd5745] <= 32'hbb4cc35d;
        mem[14'd5746] <= 32'h3bec31c8;
        mem[14'd5747] <= 32'hbc8372a2;
        mem[14'd5748] <= 32'h3c7429d9;
        mem[14'd5749] <= 32'hbd5b0e84;
        mem[14'd5750] <= 32'hbd0d43fc;
        mem[14'd5751] <= 32'hbd51dbe4;
        mem[14'd5752] <= 32'h3d1b65e7;
        mem[14'd5753] <= 32'h3b3d0e12;
        mem[14'd5754] <= 32'hbc355f9e;
        mem[14'd5755] <= 32'hbe879f7c;
        mem[14'd5756] <= 32'hbe46061f;
        mem[14'd5757] <= 32'hbe608c07;
        mem[14'd5758] <= 32'hbda92946;
        mem[14'd5759] <= 32'hbe16075a;
        mem[14'd5760] <= 32'hbe18662f;
        mem[14'd5761] <= 32'hbc5364d8;
        mem[14'd5762] <= 32'h3db24209;
        mem[14'd5763] <= 32'h3e2da38d;
        mem[14'd5764] <= 32'h3e113382;
        mem[14'd5765] <= 32'h3df4b861;
        mem[14'd5766] <= 32'h3df21b36;
        mem[14'd5767] <= 32'h3e3c59b6;
        mem[14'd5768] <= 32'h3d91d02d;
        mem[14'd5769] <= 32'hbca111c4;
        mem[14'd5770] <= 32'h3ca5865e;
        mem[14'd5771] <= 32'hbc81bb2d;
        mem[14'd5772] <= 32'h3c0b30f0;
        mem[14'd5773] <= 32'h3c1eb3da;
        mem[14'd5774] <= 32'hbc286e8f;
        mem[14'd5775] <= 32'hbc64a13b;
        mem[14'd5776] <= 32'h3c4098d9;
        mem[14'd5777] <= 32'hbdaad0db;
        mem[14'd5778] <= 32'hbdc6127e;
        mem[14'd5779] <= 32'hbd28f510;
        mem[14'd5780] <= 32'hbd530405;
        mem[14'd5781] <= 32'hbdd8af18;
        mem[14'd5782] <= 32'hbe66b85e;
        mem[14'd5783] <= 32'hbe5349e5;
        mem[14'd5784] <= 32'hbe27cc51;
        mem[14'd5785] <= 32'hbe72c7f7;
        mem[14'd5786] <= 32'hbe477480;
        mem[14'd5787] <= 32'hbe010cb4;
        mem[14'd5788] <= 32'hbe5ce5fc;
        mem[14'd5789] <= 32'hbe19a8dc;
        mem[14'd5790] <= 32'hbe382583;
        mem[14'd5791] <= 32'hbe103286;
        mem[14'd5792] <= 32'hbdd6847b;
        mem[14'd5793] <= 32'hbd813904;
        mem[14'd5794] <= 32'hbcbeedb5;
        mem[14'd5795] <= 32'h3cdc9dfe;
        mem[14'd5796] <= 32'h3cd6dea2;
        mem[14'd5797] <= 32'hbcb5121a;
        mem[14'd5798] <= 32'hbba564c9;
        mem[14'd5799] <= 32'h3c1badbb;
        mem[14'd5800] <= 32'hbb1c707e;
        mem[14'd5801] <= 32'h39905a95;
        mem[14'd5802] <= 32'hbb092a06;
        mem[14'd5803] <= 32'hbcc4aad5;
        mem[14'd5804] <= 32'hbcf29df8;
        mem[14'd5805] <= 32'hbd80a7be;
        mem[14'd5806] <= 32'hbe1f4b23;
        mem[14'd5807] <= 32'hbd9b005b;
        mem[14'd5808] <= 32'hbdb68012;
        mem[14'd5809] <= 32'hbe0f062e;
        mem[14'd5810] <= 32'hbe557a16;
        mem[14'd5811] <= 32'hbdf8d8a9;
        mem[14'd5812] <= 32'hbe23139a;
        mem[14'd5813] <= 32'hbe8791cb;
        mem[14'd5814] <= 32'hbe2a6716;
        mem[14'd5815] <= 32'hbe1ba65a;
        mem[14'd5816] <= 32'hbe927ce2;
        mem[14'd5817] <= 32'hbe6ec399;
        mem[14'd5818] <= 32'hbe9a2504;
        mem[14'd5819] <= 32'hbeaa8114;
        mem[14'd5820] <= 32'hbe829dc2;
        mem[14'd5821] <= 32'hbe4bd760;
        mem[14'd5822] <= 32'hbe564229;
        mem[14'd5823] <= 32'hbe14be06;
        mem[14'd5824] <= 32'hbc88eb11;
        mem[14'd5825] <= 32'hbd5e2c0a;
        mem[14'd5826] <= 32'hbca3f9b1;
        mem[14'd5827] <= 32'h3c2cfed8;
        mem[14'd5828] <= 32'h3b86b44d;
        mem[14'd5829] <= 32'h3c42b005;
        mem[14'd5830] <= 32'hbc29f2fb;
        mem[14'd5831] <= 32'hbc52bd1a;
        mem[14'd5832] <= 32'hbc370e5f;
        mem[14'd5833] <= 32'hbdaf9275;
        mem[14'd5834] <= 32'hbe228fcf;
        mem[14'd5835] <= 32'hbe003d16;
        mem[14'd5836] <= 32'hbde0a6ce;
        mem[14'd5837] <= 32'hbdf86f48;
        mem[14'd5838] <= 32'hbe5b1bf7;
        mem[14'd5839] <= 32'hbe0f61dc;
        mem[14'd5840] <= 32'hbe3e8624;
        mem[14'd5841] <= 32'hbe51558f;
        mem[14'd5842] <= 32'hbe8dccf0;
        mem[14'd5843] <= 32'hbeb70d70;
        mem[14'd5844] <= 32'hbebfb158;
        mem[14'd5845] <= 32'hbec81912;
        mem[14'd5846] <= 32'hbf10eec7;
        mem[14'd5847] <= 32'hbeff5b54;
        mem[14'd5848] <= 32'hbec05146;
        mem[14'd5849] <= 32'hbe92475c;
        mem[14'd5850] <= 32'hbea170b6;
        mem[14'd5851] <= 32'hbea99484;
        mem[14'd5852] <= 32'hbe69fdb3;
        mem[14'd5853] <= 32'hbe128cc8;
        mem[14'd5854] <= 32'hbd65736c;
        mem[14'd5855] <= 32'hbbb4eba5;
        mem[14'd5856] <= 32'h3a9c8b77;
        mem[14'd5857] <= 32'hbc99006d;
        mem[14'd5858] <= 32'hbb735cc0;
        mem[14'd5859] <= 32'hbd051834;
        mem[14'd5860] <= 32'hbcabd938;
        mem[14'd5861] <= 32'hbe086f53;
        mem[14'd5862] <= 32'hbe35edc9;
        mem[14'd5863] <= 32'hbd7684e5;
        mem[14'd5864] <= 32'hbd31804a;
        mem[14'd5865] <= 32'hbe3158d6;
        mem[14'd5866] <= 32'hbe5a3b1c;
        mem[14'd5867] <= 32'hbe1b29fa;
        mem[14'd5868] <= 32'hbe3ef411;
        mem[14'd5869] <= 32'hbe93fbc9;
        mem[14'd5870] <= 32'hbe6a740d;
        mem[14'd5871] <= 32'hbebe26d8;
        mem[14'd5872] <= 32'hbef551e1;
        mem[14'd5873] <= 32'hbf209398;
        mem[14'd5874] <= 32'hbf127ac5;
        mem[14'd5875] <= 32'hbef744ff;
        mem[14'd5876] <= 32'hbead9246;
        mem[14'd5877] <= 32'hbe97b0c2;
        mem[14'd5878] <= 32'hbeca7b42;
        mem[14'd5879] <= 32'hbe926097;
        mem[14'd5880] <= 32'hbe845e8d;
        mem[14'd5881] <= 32'hbe51cd55;
        mem[14'd5882] <= 32'hbda8ac72;
        mem[14'd5883] <= 32'hbc385633;
        mem[14'd5884] <= 32'hbc8894af;
        mem[14'd5885] <= 32'hbb7c7739;
        mem[14'd5886] <= 32'hbc54a100;
        mem[14'd5887] <= 32'hbcc480bc;
        mem[14'd5888] <= 32'hbd5281fc;
        mem[14'd5889] <= 32'hbdf10ffc;
        mem[14'd5890] <= 32'hbde96829;
        mem[14'd5891] <= 32'h3caf147b;
        mem[14'd5892] <= 32'h3c8f6008;
        mem[14'd5893] <= 32'hbdf23176;
        mem[14'd5894] <= 32'hbd9395e2;
        mem[14'd5895] <= 32'hbe00e089;
        mem[14'd5896] <= 32'hbe3fd3b3;
        mem[14'd5897] <= 32'hbdcd1726;
        mem[14'd5898] <= 32'hbe808881;
        mem[14'd5899] <= 32'hbee49985;
        mem[14'd5900] <= 32'hbee82342;
        mem[14'd5901] <= 32'hbee454a2;
        mem[14'd5902] <= 32'hbedac7da;
        mem[14'd5903] <= 32'hbec49095;
        mem[14'd5904] <= 32'hbe850169;
        mem[14'd5905] <= 32'hbe915775;
        mem[14'd5906] <= 32'hbe95def4;
        mem[14'd5907] <= 32'hbe13639a;
        mem[14'd5908] <= 32'hbe472098;
        mem[14'd5909] <= 32'hbe77070c;
        mem[14'd5910] <= 32'hbdc0eacd;
        mem[14'd5911] <= 32'hbc5387a2;
        mem[14'd5912] <= 32'hbafa2644;
        mem[14'd5913] <= 32'hbc3f2413;
        mem[14'd5914] <= 32'hbc1aa818;
        mem[14'd5915] <= 32'hbcff6094;
        mem[14'd5916] <= 32'hbd549d22;
        mem[14'd5917] <= 32'hbca7dfa9;
        mem[14'd5918] <= 32'hbd108018;
        mem[14'd5919] <= 32'h3de09937;
        mem[14'd5920] <= 32'h3d9c7edb;
        mem[14'd5921] <= 32'h3deb2df5;
        mem[14'd5922] <= 32'h3d33d9a6;
        mem[14'd5923] <= 32'hbd23510d;
        mem[14'd5924] <= 32'h3d8549e1;
        mem[14'd5925] <= 32'h3de2f967;
        mem[14'd5926] <= 32'hbe4bce8c;
        mem[14'd5927] <= 32'hbf0049ce;
        mem[14'd5928] <= 32'hbe8d8db6;
        mem[14'd5929] <= 32'hbea5566b;
        mem[14'd5930] <= 32'hbe8d56c9;
        mem[14'd5931] <= 32'hbe3eeb19;
        mem[14'd5932] <= 32'hbe0c999e;
        mem[14'd5933] <= 32'hbc65d64e;
        mem[14'd5934] <= 32'h3bd4195c;
        mem[14'd5935] <= 32'h3e35881f;
        mem[14'd5936] <= 32'hbcf4992e;
        mem[14'd5937] <= 32'hbe435f77;
        mem[14'd5938] <= 32'hbde085f8;
        mem[14'd5939] <= 32'hbb865ae6;
        mem[14'd5940] <= 32'h3bafea71;
        mem[14'd5941] <= 32'hbc4aaf33;
        mem[14'd5942] <= 32'h3c3f7ee3;
        mem[14'd5943] <= 32'hbccd5d79;
        mem[14'd5944] <= 32'hbda80eb4;
        mem[14'd5945] <= 32'h3aef6bfe;
        mem[14'd5946] <= 32'h3e1344ec;
        mem[14'd5947] <= 32'h3e3a76d6;
        mem[14'd5948] <= 32'h3dfd32fa;
        mem[14'd5949] <= 32'h3e13e412;
        mem[14'd5950] <= 32'h3d39d276;
        mem[14'd5951] <= 32'h3e526757;
        mem[14'd5952] <= 32'h3e46aa40;
        mem[14'd5953] <= 32'h3e0992dc;
        mem[14'd5954] <= 32'hbe657b15;
        mem[14'd5955] <= 32'hbe96e5c0;
        mem[14'd5956] <= 32'hbd96098a;
        mem[14'd5957] <= 32'hbe08b2f3;
        mem[14'd5958] <= 32'hbe2e0a78;
        mem[14'd5959] <= 32'hbe7bca1b;
        mem[14'd5960] <= 32'hbdc6c65e;
        mem[14'd5961] <= 32'h3dc602c5;
        mem[14'd5962] <= 32'h3e8be28f;
        mem[14'd5963] <= 32'h3ef6f2bd;
        mem[14'd5964] <= 32'h3e55645c;
        mem[14'd5965] <= 32'hbe068258;
        mem[14'd5966] <= 32'hbdbc3c77;
        mem[14'd5967] <= 32'hbc5721b0;
        mem[14'd5968] <= 32'hbbbe315b;
        mem[14'd5969] <= 32'hbc881323;
        mem[14'd5970] <= 32'hbb449247;
        mem[14'd5971] <= 32'hbd192d23;
        mem[14'd5972] <= 32'hbdaca3bc;
        mem[14'd5973] <= 32'h3dbac158;
        mem[14'd5974] <= 32'h3e859a82;
        mem[14'd5975] <= 32'h3db6ef11;
        mem[14'd5976] <= 32'h3dc874a5;
        mem[14'd5977] <= 32'h3df86360;
        mem[14'd5978] <= 32'h3e2d0485;
        mem[14'd5979] <= 32'h3dfc5df2;
        mem[14'd5980] <= 32'h3e216258;
        mem[14'd5981] <= 32'h3cf388f4;
        mem[14'd5982] <= 32'hbe128702;
        mem[14'd5983] <= 32'h3d4722dc;
        mem[14'd5984] <= 32'h3ccc6b37;
        mem[14'd5985] <= 32'hbe2c281a;
        mem[14'd5986] <= 32'hbe2508da;
        mem[14'd5987] <= 32'hbcc01c98;
        mem[14'd5988] <= 32'hbd8e9139;
        mem[14'd5989] <= 32'h3e09293f;
        mem[14'd5990] <= 32'h3eb4b50b;
        mem[14'd5991] <= 32'h3f0ff317;
        mem[14'd5992] <= 32'h3e8dad80;
        mem[14'd5993] <= 32'hbde7a543;
        mem[14'd5994] <= 32'hbde058ee;
        mem[14'd5995] <= 32'hbcb5c77e;
        mem[14'd5996] <= 32'h3b4f4f57;
        mem[14'd5997] <= 32'hbc837da2;
        mem[14'd5998] <= 32'hbc4aacf1;
        mem[14'd5999] <= 32'hbc53f14e;
        mem[14'd6000] <= 32'hbe114dc4;
        mem[14'd6001] <= 32'h3d906b76;
        mem[14'd6002] <= 32'h3e4b3c19;
        mem[14'd6003] <= 32'h3df9c0ef;
        mem[14'd6004] <= 32'h3e230a9f;
        mem[14'd6005] <= 32'h3e52c022;
        mem[14'd6006] <= 32'h3e78f5a1;
        mem[14'd6007] <= 32'h3eb6f867;
        mem[14'd6008] <= 32'h3e197417;
        mem[14'd6009] <= 32'hbd39b289;
        mem[14'd6010] <= 32'hbcabb36c;
        mem[14'd6011] <= 32'h3dc4e9a3;
        mem[14'd6012] <= 32'h3da4e89a;
        mem[14'd6013] <= 32'hbe5a042a;
        mem[14'd6014] <= 32'hbe2bec91;
        mem[14'd6015] <= 32'hbd19b1ff;
        mem[14'd6016] <= 32'h3c8465df;
        mem[14'd6017] <= 32'h3e0e2d09;
        mem[14'd6018] <= 32'h3ea5a167;
        mem[14'd6019] <= 32'h3ed048ae;
        mem[14'd6020] <= 32'h3e44d0f3;
        mem[14'd6021] <= 32'hbd83b916;
        mem[14'd6022] <= 32'hbdd31a37;
        mem[14'd6023] <= 32'h39f72356;
        mem[14'd6024] <= 32'hbbe9ee21;
        mem[14'd6025] <= 32'h3b7b9add;
        mem[14'd6026] <= 32'hb9d36a1b;
        mem[14'd6027] <= 32'hbd570157;
        mem[14'd6028] <= 32'hbe5dced5;
        mem[14'd6029] <= 32'h3c4bffca;
        mem[14'd6030] <= 32'h3e51d533;
        mem[14'd6031] <= 32'h3e5cef9e;
        mem[14'd6032] <= 32'h3e57a909;
        mem[14'd6033] <= 32'h3e349838;
        mem[14'd6034] <= 32'h3e95405b;
        mem[14'd6035] <= 32'h3ebaa412;
        mem[14'd6036] <= 32'h3e2ad986;
        mem[14'd6037] <= 32'h3d6c6f0f;
        mem[14'd6038] <= 32'h3e422a1a;
        mem[14'd6039] <= 32'h3de50a23;
        mem[14'd6040] <= 32'hbb9c2f63;
        mem[14'd6041] <= 32'hbd9df337;
        mem[14'd6042] <= 32'hbdbccf27;
        mem[14'd6043] <= 32'hbc0c9480;
        mem[14'd6044] <= 32'h3df59f41;
        mem[14'd6045] <= 32'h3e04d58e;
        mem[14'd6046] <= 32'h3ddc9029;
        mem[14'd6047] <= 32'h3e5866be;
        mem[14'd6048] <= 32'h3db9269b;
        mem[14'd6049] <= 32'hbd5cf69c;
        mem[14'd6050] <= 32'hbdc9111d;
        mem[14'd6051] <= 32'hbd0faeae;
        mem[14'd6052] <= 32'hbbec788a;
        mem[14'd6053] <= 32'hbaffee0f;
        mem[14'd6054] <= 32'h3b0a553a;
        mem[14'd6055] <= 32'hbda3b7d1;
        mem[14'd6056] <= 32'hbe6a1653;
        mem[14'd6057] <= 32'h3b7a399b;
        mem[14'd6058] <= 32'h3e5d48d1;
        mem[14'd6059] <= 32'h3e8f6a18;
        mem[14'd6060] <= 32'h3e78a395;
        mem[14'd6061] <= 32'h3e97d7d9;
        mem[14'd6062] <= 32'h3ec76ecd;
        mem[14'd6063] <= 32'h3f0b8957;
        mem[14'd6064] <= 32'h3d91ac26;
        mem[14'd6065] <= 32'h3cfa2549;
        mem[14'd6066] <= 32'h3e332c16;
        mem[14'd6067] <= 32'h3d8875e0;
        mem[14'd6068] <= 32'hbd97501e;
        mem[14'd6069] <= 32'hbe25ec48;
        mem[14'd6070] <= 32'h3da854cc;
        mem[14'd6071] <= 32'h3deeec40;
        mem[14'd6072] <= 32'h3c24f86c;
        mem[14'd6073] <= 32'h3b256d42;
        mem[14'd6074] <= 32'hbc915c32;
        mem[14'd6075] <= 32'h3d8beea7;
        mem[14'd6076] <= 32'h3d0c5fe5;
        mem[14'd6077] <= 32'hbd9ce8bf;
        mem[14'd6078] <= 32'hbdba8171;
        mem[14'd6079] <= 32'hbc4968f9;
        mem[14'd6080] <= 32'hba2f2df3;
        mem[14'd6081] <= 32'h3bf41d73;
        mem[14'd6082] <= 32'h3c7c9fd3;
        mem[14'd6083] <= 32'hbd9c388c;
        mem[14'd6084] <= 32'hbe90d66b;
        mem[14'd6085] <= 32'hbdf1dddc;
        mem[14'd6086] <= 32'h3dd855f4;
        mem[14'd6087] <= 32'h3e7430a3;
        mem[14'd6088] <= 32'h3e8ba20c;
        mem[14'd6089] <= 32'h3e936efc;
        mem[14'd6090] <= 32'h3efe6c7a;
        mem[14'd6091] <= 32'h3efcc98c;
        mem[14'd6092] <= 32'h3e2d8918;
        mem[14'd6093] <= 32'h3dd32f8b;
        mem[14'd6094] <= 32'h3e0c31d2;
        mem[14'd6095] <= 32'hbc0588c3;
        mem[14'd6096] <= 32'hbd9243f4;
        mem[14'd6097] <= 32'h3d3d30fe;
        mem[14'd6098] <= 32'h3e195632;
        mem[14'd6099] <= 32'h3e0ee9f7;
        mem[14'd6100] <= 32'h3d2db4c1;
        mem[14'd6101] <= 32'h3c5dd285;
        mem[14'd6102] <= 32'h3d5d3e84;
        mem[14'd6103] <= 32'h3d29d932;
        mem[14'd6104] <= 32'hbcbe8b91;
        mem[14'd6105] <= 32'hbd1bd097;
        mem[14'd6106] <= 32'hbd3c2afd;
        mem[14'd6107] <= 32'h3a3420d8;
        mem[14'd6108] <= 32'hbc329cd9;
        mem[14'd6109] <= 32'h3c2a99ef;
        mem[14'd6110] <= 32'hbc009a50;
        mem[14'd6111] <= 32'hbda07ad5;
        mem[14'd6112] <= 32'hbe6f9590;
        mem[14'd6113] <= 32'hbe6c76b1;
        mem[14'd6114] <= 32'hbd185f48;
        mem[14'd6115] <= 32'h3e3acd66;
        mem[14'd6116] <= 32'h3e45f39c;
        mem[14'd6117] <= 32'h3e84b69c;
        mem[14'd6118] <= 32'h3e950188;
        mem[14'd6119] <= 32'h3eadb534;
        mem[14'd6120] <= 32'h3f007a60;
        mem[14'd6121] <= 32'h3e825569;
        mem[14'd6122] <= 32'h3d8672a1;
        mem[14'd6123] <= 32'h3d8b166a;
        mem[14'd6124] <= 32'h3e4c2c01;
        mem[14'd6125] <= 32'h3e6c395c;
        mem[14'd6126] <= 32'h3e7b6117;
        mem[14'd6127] <= 32'h3d37ae55;
        mem[14'd6128] <= 32'h3cb61907;
        mem[14'd6129] <= 32'h3d67e85e;
        mem[14'd6130] <= 32'h3c9a5d4f;
        mem[14'd6131] <= 32'h3d1928c6;
        mem[14'd6132] <= 32'hbd3b96ef;
        mem[14'd6133] <= 32'hbca0f002;
        mem[14'd6134] <= 32'hbcedcce9;
        mem[14'd6135] <= 32'hbc90fd5b;
        mem[14'd6136] <= 32'h3b92e369;
        mem[14'd6137] <= 32'h3b012f8c;
        mem[14'd6138] <= 32'hbc8e212e;
        mem[14'd6139] <= 32'hbd88814b;
        mem[14'd6140] <= 32'hbe42f416;
        mem[14'd6141] <= 32'hbe65f577;
        mem[14'd6142] <= 32'hbda96cbd;
        mem[14'd6143] <= 32'h3d59c575;
        mem[14'd6144] <= 32'h3d69e8d9;
        mem[14'd6145] <= 32'h3e708513;
        mem[14'd6146] <= 32'h3eb141c3;
        mem[14'd6147] <= 32'h3f0b6a35;
        mem[14'd6148] <= 32'h3f0964c3;
        mem[14'd6149] <= 32'h3e813950;
        mem[14'd6150] <= 32'h3e8cc775;
        mem[14'd6151] <= 32'h3e6f917a;
        mem[14'd6152] <= 32'h3e6a69c0;
        mem[14'd6153] <= 32'h3e30d5bc;
        mem[14'd6154] <= 32'h3da99d5e;
        mem[14'd6155] <= 32'h3d99894b;
        mem[14'd6156] <= 32'h3d997396;
        mem[14'd6157] <= 32'h3dadb0fd;
        mem[14'd6158] <= 32'h3dad40bf;
        mem[14'd6159] <= 32'hbc381874;
        mem[14'd6160] <= 32'hbd882380;
        mem[14'd6161] <= 32'hbdb31651;
        mem[14'd6162] <= 32'hbd246cbb;
        mem[14'd6163] <= 32'hbc2170fd;
        mem[14'd6164] <= 32'hbb3663d2;
        mem[14'd6165] <= 32'hbc0d88fc;
        mem[14'd6166] <= 32'h3b348ff1;
        mem[14'd6167] <= 32'hbd2b9a06;
        mem[14'd6168] <= 32'hbe1ae537;
        mem[14'd6169] <= 32'hbe7d738e;
        mem[14'd6170] <= 32'hbe35ea45;
        mem[14'd6171] <= 32'h3d09ffae;
        mem[14'd6172] <= 32'h3c950b54;
        mem[14'd6173] <= 32'h3e560c15;
        mem[14'd6174] <= 32'h3ebedacc;
        mem[14'd6175] <= 32'h3ea28f92;
        mem[14'd6176] <= 32'h3ee698a4;
        mem[14'd6177] <= 32'h3eb27d1f;
        mem[14'd6178] <= 32'h3f03a6ef;
        mem[14'd6179] <= 32'h3eb41af4;
        mem[14'd6180] <= 32'h3e4e8502;
        mem[14'd6181] <= 32'h3dba7068;
        mem[14'd6182] <= 32'h3e541262;
        mem[14'd6183] <= 32'h3dcdaae6;
        mem[14'd6184] <= 32'h3dd88614;
        mem[14'd6185] <= 32'h3cce0bb0;
        mem[14'd6186] <= 32'hbdb1b35e;
        mem[14'd6187] <= 32'hbd0c7c3b;
        mem[14'd6188] <= 32'hbda345ec;
        mem[14'd6189] <= 32'hbd43326b;
        mem[14'd6190] <= 32'h3b9fb661;
        mem[14'd6191] <= 32'hbb5d94c9;
        mem[14'd6192] <= 32'h3bc619cd;
        mem[14'd6193] <= 32'h3c4623b3;
        mem[14'd6194] <= 32'h3c0f76a1;
        mem[14'd6195] <= 32'hbccea5eb;
        mem[14'd6196] <= 32'hbde5e214;
        mem[14'd6197] <= 32'hbe651d4f;
        mem[14'd6198] <= 32'hbe9db9e1;
        mem[14'd6199] <= 32'hbdb449a1;
        mem[14'd6200] <= 32'h3de47c60;
        mem[14'd6201] <= 32'h3e430890;
        mem[14'd6202] <= 32'h3e8219dc;
        mem[14'd6203] <= 32'h3ea5335b;
        mem[14'd6204] <= 32'h3f02d70c;
        mem[14'd6205] <= 32'h3f034aac;
        mem[14'd6206] <= 32'h3ee6f93f;
        mem[14'd6207] <= 32'h3e8b024c;
        mem[14'd6208] <= 32'h3e66c1e7;
        mem[14'd6209] <= 32'h3e8dde16;
        mem[14'd6210] <= 32'h3e89b921;
        mem[14'd6211] <= 32'h3dc9456c;
        mem[14'd6212] <= 32'h3ceeb371;
        mem[14'd6213] <= 32'hbd957bac;
        mem[14'd6214] <= 32'hbd29d5cc;
        mem[14'd6215] <= 32'hbd3631a4;
        mem[14'd6216] <= 32'hbd05393c;
        mem[14'd6217] <= 32'hbd16d734;
        mem[14'd6218] <= 32'hbb701c27;
        mem[14'd6219] <= 32'hbc6ef8a2;
        mem[14'd6220] <= 32'h3a18632e;
        mem[14'd6221] <= 32'hbbaedd2e;
        mem[14'd6222] <= 32'h3c606da3;
        mem[14'd6223] <= 32'hbb356aa0;
        mem[14'd6224] <= 32'hbd33af25;
        mem[14'd6225] <= 32'hbe0b89a7;
        mem[14'd6226] <= 32'hbe8a19fe;
        mem[14'd6227] <= 32'hbe80d1b4;
        mem[14'd6228] <= 32'hbe00ce6e;
        mem[14'd6229] <= 32'hbd140f1c;
        mem[14'd6230] <= 32'h3dc0abac;
        mem[14'd6231] <= 32'h3d1c15dd;
        mem[14'd6232] <= 32'h3e4fae98;
        mem[14'd6233] <= 32'h3e291e91;
        mem[14'd6234] <= 32'h3d6208be;
        mem[14'd6235] <= 32'h3e5a0801;
        mem[14'd6236] <= 32'h3dc21820;
        mem[14'd6237] <= 32'h3d12aad5;
        mem[14'd6238] <= 32'hbd49bd75;
        mem[14'd6239] <= 32'hbd234936;
        mem[14'd6240] <= 32'hbcec35bd;
        mem[14'd6241] <= 32'hbd4d89de;
        mem[14'd6242] <= 32'hbdbeb8ce;
        mem[14'd6243] <= 32'hbdb32b42;
        mem[14'd6244] <= 32'hbd1ff65e;
        mem[14'd6245] <= 32'h3b6ba933;
        mem[14'd6246] <= 32'hbb90c309;
        mem[14'd6247] <= 32'hbc74df96;
        mem[14'd6248] <= 32'hbb4b19a4;
        mem[14'd6249] <= 32'hbc900d22;
        mem[14'd6250] <= 32'h3b742679;
        mem[14'd6251] <= 32'hbc720774;
        mem[14'd6252] <= 32'hbcb9cc3f;
        mem[14'd6253] <= 32'hbd63046f;
        mem[14'd6254] <= 32'hbdcb4e73;
        mem[14'd6255] <= 32'hbe585da4;
        mem[14'd6256] <= 32'hbe82b9b7;
        mem[14'd6257] <= 32'hbe8baaa6;
        mem[14'd6258] <= 32'hbeac2f0b;
        mem[14'd6259] <= 32'hbe9d33b3;
        mem[14'd6260] <= 32'hbe2f7a16;
        mem[14'd6261] <= 32'hbda48b41;
        mem[14'd6262] <= 32'hbda046e1;
        mem[14'd6263] <= 32'hbd8febc2;
        mem[14'd6264] <= 32'hbde0ad69;
        mem[14'd6265] <= 32'hbe11b575;
        mem[14'd6266] <= 32'hbd70d03b;
        mem[14'd6267] <= 32'hbd00d0f1;
        mem[14'd6268] <= 32'hbcef53d2;
        mem[14'd6269] <= 32'hbd74dd17;
        mem[14'd6270] <= 32'hbd57ec2f;
        mem[14'd6271] <= 32'hbd092087;
        mem[14'd6272] <= 32'hbc25ade1;
        mem[14'd6273] <= 32'hbc019787;
        mem[14'd6274] <= 32'hbb8a213d;
        mem[14'd6275] <= 32'h3cb57db5;
        mem[14'd6276] <= 32'hbaa2b7a7;
        mem[14'd6277] <= 32'hbc63d74e;
        mem[14'd6278] <= 32'hbc567e01;
        mem[14'd6279] <= 32'h3bfe9361;
        mem[14'd6280] <= 32'hbaf561d6;
        mem[14'd6281] <= 32'hbb211758;
        mem[14'd6282] <= 32'hbbf624c8;
        mem[14'd6283] <= 32'hbd8222db;
        mem[14'd6284] <= 32'hbdee590b;
        mem[14'd6285] <= 32'hbe246d6d;
        mem[14'd6286] <= 32'hbe594344;
        mem[14'd6287] <= 32'hbe9077de;
        mem[14'd6288] <= 32'hbe8e94eb;
        mem[14'd6289] <= 32'hbe93c0a1;
        mem[14'd6290] <= 32'hbe8b07e1;
        mem[14'd6291] <= 32'hbe73f759;
        mem[14'd6292] <= 32'hbe231428;
        mem[14'd6293] <= 32'hbde268c6;
        mem[14'd6294] <= 32'hbdb6677c;
        mem[14'd6295] <= 32'hbd89662e;
        mem[14'd6296] <= 32'hbd3af074;
        mem[14'd6297] <= 32'hbd4219a4;
        mem[14'd6298] <= 32'hbd4015b9;
        mem[14'd6299] <= 32'h3c06839b;
        mem[14'd6300] <= 32'hbb9bb6b0;
        mem[14'd6301] <= 32'h3c5fe84b;
        mem[14'd6302] <= 32'h3bb46288;
        mem[14'd6303] <= 32'hbbba19ea;
        mem[14'd6304] <= 32'hbb8d8cc2;
        mem[14'd6305] <= 32'h3c477274;
        mem[14'd6306] <= 32'h3c21038a;
        mem[14'd6307] <= 32'h3bb62642;
        mem[14'd6308] <= 32'h3c61d02b;
        mem[14'd6309] <= 32'h3c024d7f;
        mem[14'd6310] <= 32'h3b286906;
        mem[14'd6311] <= 32'hbcbf5359;
        mem[14'd6312] <= 32'hbcae841d;
        mem[14'd6313] <= 32'hbd63f780;
        mem[14'd6314] <= 32'hbd0a11f8;
        mem[14'd6315] <= 32'hbd02eaa5;
        mem[14'd6316] <= 32'hbd4a6cc4;
        mem[14'd6317] <= 32'hbd989779;
        mem[14'd6318] <= 32'hbd9ffbd5;
        mem[14'd6319] <= 32'hbda31a80;
        mem[14'd6320] <= 32'hbd84532e;
        mem[14'd6321] <= 32'hbd415973;
        mem[14'd6322] <= 32'hbc8edea3;
        mem[14'd6323] <= 32'hbc9aad51;
        mem[14'd6324] <= 32'hbcc3aaaa;
        mem[14'd6325] <= 32'hbc96b5f8;
        mem[14'd6326] <= 32'h3c293b49;
        mem[14'd6327] <= 32'hbb83df97;
        mem[14'd6328] <= 32'hbc49b1d2;
        mem[14'd6329] <= 32'hbb5494df;
        mem[14'd6330] <= 32'h39e1f751;
        mem[14'd6331] <= 32'h3bf7ca50;
        mem[14'd6332] <= 32'hbbeff22b;
        mem[14'd6333] <= 32'hbb137367;
        mem[14'd6334] <= 32'h3c14e629;
        mem[14'd6335] <= 32'h3ca3c384;
        mem[14'd6336] <= 32'hbc8fef1a;
        mem[14'd6337] <= 32'hbbe7d233;
        mem[14'd6338] <= 32'hba302ec6;
        mem[14'd6339] <= 32'h3c219a90;
        mem[14'd6340] <= 32'hbc0464db;
        mem[14'd6341] <= 32'hbb9c62a8;
        mem[14'd6342] <= 32'hbb4c6a32;
        mem[14'd6343] <= 32'hbc3f67a7;
        mem[14'd6344] <= 32'hbc58c7ee;
        mem[14'd6345] <= 32'hbca470d6;
        mem[14'd6346] <= 32'hb98cec4a;
        mem[14'd6347] <= 32'hbb69e6aa;
        mem[14'd6348] <= 32'hbca548e2;
        mem[14'd6349] <= 32'hbba30d6a;
        mem[14'd6350] <= 32'h3b69ca11;
        mem[14'd6351] <= 32'hbc94d24c;
        mem[14'd6352] <= 32'h3c69c793;
        mem[14'd6353] <= 32'h3b90d4bf;
        mem[14'd6354] <= 32'h3ba3b7e9;
        mem[14'd6355] <= 32'h3b1bddd6;
        mem[14'd6356] <= 32'h3bb7effd;
        mem[14'd6357] <= 32'hbbdafe09;
        mem[14'd6358] <= 32'hbc020d5f;
        mem[14'd6359] <= 32'hbb9a76eb;
        mem[14'd6360] <= 32'h3ca86201;
        mem[14'd6361] <= 32'hbcce5ddd;
        mem[14'd6362] <= 32'h3b8d7b19;
        mem[14'd6363] <= 32'hbb916ccb;
        mem[14'd6364] <= 32'h3babd4a3;
        mem[14'd6365] <= 32'h3b805cb1;
        mem[14'd6366] <= 32'hbbfcb4d4;
        mem[14'd6367] <= 32'hbc950309;
        mem[14'd6368] <= 32'hbbe3d150;
        mem[14'd6369] <= 32'h3ba5f4de;
        mem[14'd6370] <= 32'hbb4c4ea3;
        mem[14'd6371] <= 32'h3c0b7d81;
        mem[14'd6372] <= 32'hba009063;
        mem[14'd6373] <= 32'h3c8a8765;
        mem[14'd6374] <= 32'hbc1b8a70;
        mem[14'd6375] <= 32'hbb9f72bc;
        mem[14'd6376] <= 32'h3bdc72b4;
        mem[14'd6377] <= 32'hbcefa08c;
        mem[14'd6378] <= 32'h3c46161f;
        mem[14'd6379] <= 32'h3b824098;
        mem[14'd6380] <= 32'h3b839ff1;
        mem[14'd6381] <= 32'hbaaffe68;
        mem[14'd6382] <= 32'h3c97e329;
        mem[14'd6383] <= 32'h3afc9c1e;
        mem[14'd6384] <= 32'hbbef4738;
        mem[14'd6385] <= 32'h3ba37321;
        mem[14'd6386] <= 32'h3b0e68b1;
        mem[14'd6387] <= 32'hbb13b0b9;
        mem[14'd6388] <= 32'hbc54b6a2;
        mem[14'd6389] <= 32'hb94f6abc;
        mem[14'd6390] <= 32'h3b74e025;
        mem[14'd6391] <= 32'h3bfea865;
        mem[14'd6392] <= 32'h3c8ebd0f;
        mem[14'd6393] <= 32'h3c4ed450;
        mem[14'd6394] <= 32'hbbb3638f;
        mem[14'd6395] <= 32'hb8919f9e;
        mem[14'd6396] <= 32'h3c36196e;
        mem[14'd6397] <= 32'hbc3174f4;
        mem[14'd6398] <= 32'hbc59a36f;
        mem[14'd6399] <= 32'h3b821315;
        mem[14'd6400] <= 32'hbc29d8d3;
        mem[14'd6401] <= 32'hbb19f6dc;
        mem[14'd6402] <= 32'hbc49095b;
        mem[14'd6403] <= 32'hbcdd7dc2;
        mem[14'd6404] <= 32'h3a75b65c;
        mem[14'd6405] <= 32'h3b764d12;
        mem[14'd6406] <= 32'hbc882b04;
        mem[14'd6407] <= 32'hbbfab520;
        mem[14'd6408] <= 32'hbb5e6350;
        mem[14'd6409] <= 32'h3c3aa8e5;
        mem[14'd6410] <= 32'hbc0dd5ef;
        mem[14'd6411] <= 32'h3b979255;
        mem[14'd6412] <= 32'h3bf41c57;
        mem[14'd6413] <= 32'hbb11e375;
        mem[14'd6414] <= 32'hbc47e2b8;
        mem[14'd6415] <= 32'hbc83e7a4;
        mem[14'd6416] <= 32'hbb80112d;
        mem[14'd6417] <= 32'hbc38c6ca;
        mem[14'd6418] <= 32'h3944a247;
        mem[14'd6419] <= 32'h3bea31af;
        mem[14'd6420] <= 32'h38bcafac;
        mem[14'd6421] <= 32'h3c7d9a92;
        mem[14'd6422] <= 32'h3c262399;
        mem[14'd6423] <= 32'h3cad7b3c;
        mem[14'd6424] <= 32'h3b534138;
        mem[14'd6425] <= 32'hbb269116;
        mem[14'd6426] <= 32'h3c299aed;
        mem[14'd6427] <= 32'h3b925f37;
        mem[14'd6428] <= 32'hbc98a867;
        mem[14'd6429] <= 32'hba723d0e;
        mem[14'd6430] <= 32'h3bbeb79e;
        mem[14'd6431] <= 32'hbbeba2a3;
        mem[14'd6432] <= 32'hbc356008;
        mem[14'd6433] <= 32'hbb866789;
        mem[14'd6434] <= 32'hbb172ea9;
        mem[14'd6435] <= 32'hbba75239;
        mem[14'd6436] <= 32'h3c38bf18;
        mem[14'd6437] <= 32'hbc130fae;
        mem[14'd6438] <= 32'h3c23df80;
        mem[14'd6439] <= 32'hbc5b0cbe;
        mem[14'd6440] <= 32'hbab83a09;
        mem[14'd6441] <= 32'hbb8c02de;
        mem[14'd6442] <= 32'h3bf78423;
        mem[14'd6443] <= 32'hbc5988c2;
        mem[14'd6444] <= 32'hbc3e482d;
        mem[14'd6445] <= 32'hbbd75c90;
        mem[14'd6446] <= 32'hbb659dc3;
        mem[14'd6447] <= 32'h3b9bcd32;
        mem[14'd6448] <= 32'h3c0a2292;
        mem[14'd6449] <= 32'h3bd6d952;
        mem[14'd6450] <= 32'hbc892cbf;
        mem[14'd6451] <= 32'h3c7466a7;
        mem[14'd6452] <= 32'hbcab5160;
        mem[14'd6453] <= 32'hbbc338eb;
        mem[14'd6454] <= 32'hbca6673e;
        mem[14'd6455] <= 32'hbd001a5e;
        mem[14'd6456] <= 32'hbc5936c5;
        mem[14'd6457] <= 32'hbbc2eaa6;
        mem[14'd6458] <= 32'hbd19e0b5;
        mem[14'd6459] <= 32'hbcb1d047;
        mem[14'd6460] <= 32'hbbfed6e3;
        mem[14'd6461] <= 32'h39eb964e;
        mem[14'd6462] <= 32'h3a6f45aa;
        mem[14'd6463] <= 32'h3b9e104e;
        mem[14'd6464] <= 32'h3b893baa;
        mem[14'd6465] <= 32'hbb921e4e;
        mem[14'd6466] <= 32'hba7315ac;
        mem[14'd6467] <= 32'h3beb96d3;
        mem[14'd6468] <= 32'h3bd9ff8d;
        mem[14'd6469] <= 32'h3c1b4f7b;
        mem[14'd6470] <= 32'h3cc7822e;
        mem[14'd6471] <= 32'h3c59773e;
        mem[14'd6472] <= 32'hbb08579f;
        mem[14'd6473] <= 32'h3bff64c6;
        mem[14'd6474] <= 32'h3c31c100;
        mem[14'd6475] <= 32'h3c2a2517;
        mem[14'd6476] <= 32'h3be9e594;
        mem[14'd6477] <= 32'h3b7cb468;
        mem[14'd6478] <= 32'h3bd19459;
        mem[14'd6479] <= 32'hbc77cd13;
        mem[14'd6480] <= 32'hbd01b0b3;
        mem[14'd6481] <= 32'hbd38575e;
        mem[14'd6482] <= 32'hbd84f696;
        mem[14'd6483] <= 32'hbdad4e85;
        mem[14'd6484] <= 32'hbd9283fd;
        mem[14'd6485] <= 32'hbd92ec05;
        mem[14'd6486] <= 32'hbd9e605c;
        mem[14'd6487] <= 32'hbd6f1150;
        mem[14'd6488] <= 32'hbd5785ed;
        mem[14'd6489] <= 32'hbd593cb3;
        mem[14'd6490] <= 32'hbd0a177d;
        mem[14'd6491] <= 32'hbcbd22ee;
        mem[14'd6492] <= 32'hbc3e9006;
        mem[14'd6493] <= 32'hbc587666;
        mem[14'd6494] <= 32'h3bc2b2ab;
        mem[14'd6495] <= 32'h3b19f810;
        mem[14'd6496] <= 32'hbbc8ded3;
        mem[14'd6497] <= 32'h3c8c1062;
        mem[14'd6498] <= 32'h3c738ab7;
        mem[14'd6499] <= 32'hbbbf3b8b;
        mem[14'd6500] <= 32'h3c7efaa9;
        mem[14'd6501] <= 32'h3c92b6a0;
        mem[14'd6502] <= 32'h3bc9e70b;
        mem[14'd6503] <= 32'h3a88f494;
        mem[14'd6504] <= 32'hbca6f5f4;
        mem[14'd6505] <= 32'hbbda91c3;
        mem[14'd6506] <= 32'h399d5f5b;
        mem[14'd6507] <= 32'hbcee45bc;
        mem[14'd6508] <= 32'hbd7d60ae;
        mem[14'd6509] <= 32'hbda80ca2;
        mem[14'd6510] <= 32'hbe2650db;
        mem[14'd6511] <= 32'hbe41ae96;
        mem[14'd6512] <= 32'hbe4c61b2;
        mem[14'd6513] <= 32'hbe59bc92;
        mem[14'd6514] <= 32'hbe7acfed;
        mem[14'd6515] <= 32'hbe6bc3ab;
        mem[14'd6516] <= 32'hbe6fac22;
        mem[14'd6517] <= 32'hbe42cdde;
        mem[14'd6518] <= 32'hbe19b0c2;
        mem[14'd6519] <= 32'hbde8b30b;
        mem[14'd6520] <= 32'hbd80d3ec;
        mem[14'd6521] <= 32'hbd8aba5a;
        mem[14'd6522] <= 32'hbc934e64;
        mem[14'd6523] <= 32'hbcf4a577;
        mem[14'd6524] <= 32'h3b32b0e5;
        mem[14'd6525] <= 32'h3b2c709f;
        mem[14'd6526] <= 32'h3bbe0fa5;
        mem[14'd6527] <= 32'hbc06e330;
        mem[14'd6528] <= 32'hbbd3892f;
        mem[14'd6529] <= 32'h3bd0ff59;
        mem[14'd6530] <= 32'h3abe7176;
        mem[14'd6531] <= 32'h3c79fecd;
        mem[14'd6532] <= 32'hbb020b1b;
        mem[14'd6533] <= 32'h3d06f854;
        mem[14'd6534] <= 32'h3cccd2bb;
        mem[14'd6535] <= 32'h3ce6d853;
        mem[14'd6536] <= 32'h3d161cba;
        mem[14'd6537] <= 32'h3c062386;
        mem[14'd6538] <= 32'hbdbaa5bf;
        mem[14'd6539] <= 32'hbe36da39;
        mem[14'd6540] <= 32'hbe4b7f8e;
        mem[14'd6541] <= 32'hbe768779;
        mem[14'd6542] <= 32'hbe9a7c71;
        mem[14'd6543] <= 32'hbea7dba6;
        mem[14'd6544] <= 32'hbeaf6904;
        mem[14'd6545] <= 32'hbecfd4a2;
        mem[14'd6546] <= 32'hbec07563;
        mem[14'd6547] <= 32'hbeb40b3d;
        mem[14'd6548] <= 32'hbe9f1200;
        mem[14'd6549] <= 32'hbe4a0e9c;
        mem[14'd6550] <= 32'hbe066fa5;
        mem[14'd6551] <= 32'hbd7d1ac4;
        mem[14'd6552] <= 32'hbc70c416;
        mem[14'd6553] <= 32'hbc061041;
        mem[14'd6554] <= 32'hbc08c063;
        mem[14'd6555] <= 32'hbbd8d9f2;
        mem[14'd6556] <= 32'h3bda377b;
        mem[14'd6557] <= 32'hbcb75572;
        mem[14'd6558] <= 32'h3ba4acf0;
        mem[14'd6559] <= 32'h3d3a76de;
        mem[14'd6560] <= 32'h3c3dbf92;
        mem[14'd6561] <= 32'h3dcb73e2;
        mem[14'd6562] <= 32'h3e15553c;
        mem[14'd6563] <= 32'h3e1df767;
        mem[14'd6564] <= 32'h3e4223b8;
        mem[14'd6565] <= 32'h3df22c32;
        mem[14'd6566] <= 32'h3e32b63a;
        mem[14'd6567] <= 32'h3e6a27f2;
        mem[14'd6568] <= 32'h3dd40d36;
        mem[14'd6569] <= 32'hbdbe88ac;
        mem[14'd6570] <= 32'hbd9e9654;
        mem[14'd6571] <= 32'hbcb8f468;
        mem[14'd6572] <= 32'hbc358881;
        mem[14'd6573] <= 32'h3bf9a413;
        mem[14'd6574] <= 32'hbdc73c10;
        mem[14'd6575] <= 32'hbde9e113;
        mem[14'd6576] <= 32'hbe0113cc;
        mem[14'd6577] <= 32'hbd908397;
        mem[14'd6578] <= 32'hbdcc78f9;
        mem[14'd6579] <= 32'hbdfbaa23;
        mem[14'd6580] <= 32'hbd6e24bc;
        mem[14'd6581] <= 32'hbd24605e;
        mem[14'd6582] <= 32'hba50c1f8;
        mem[14'd6583] <= 32'h3c006b5c;
        mem[14'd6584] <= 32'hbb3e4aba;
        mem[14'd6585] <= 32'h3c3a6de0;
        mem[14'd6586] <= 32'h3c93b9b1;
        mem[14'd6587] <= 32'h3ded54ad;
        mem[14'd6588] <= 32'h3d9b850e;
        mem[14'd6589] <= 32'h3df6119e;
        mem[14'd6590] <= 32'h3e62ba0a;
        mem[14'd6591] <= 32'h3e928eb1;
        mem[14'd6592] <= 32'h3e15179e;
        mem[14'd6593] <= 32'h3e67ab54;
        mem[14'd6594] <= 32'h3e8a2e4f;
        mem[14'd6595] <= 32'h3e6d7828;
        mem[14'd6596] <= 32'h3e4f26b2;
        mem[14'd6597] <= 32'h3dfb3b69;
        mem[14'd6598] <= 32'hbd40f4ac;
        mem[14'd6599] <= 32'h3dc18b69;
        mem[14'd6600] <= 32'h3e514e5d;
        mem[14'd6601] <= 32'h3e9448ad;
        mem[14'd6602] <= 32'h3e99044a;
        mem[14'd6603] <= 32'h3e123267;
        mem[14'd6604] <= 32'h3e2f183f;
        mem[14'd6605] <= 32'h3d7dc9d7;
        mem[14'd6606] <= 32'h3c95f3f1;
        mem[14'd6607] <= 32'hbd09d0e0;
        mem[14'd6608] <= 32'hbdaca804;
        mem[14'd6609] <= 32'hbd249b07;
        mem[14'd6610] <= 32'hbb9c2521;
        mem[14'd6611] <= 32'h3cae1ce9;
        mem[14'd6612] <= 32'h3c8aa723;
        mem[14'd6613] <= 32'h3ba43d4c;
        mem[14'd6614] <= 32'h3d7ec2a2;
        mem[14'd6615] <= 32'h3e335cf8;
        mem[14'd6616] <= 32'h3e43a6fb;
        mem[14'd6617] <= 32'h3e5a36b3;
        mem[14'd6618] <= 32'h3e752197;
        mem[14'd6619] <= 32'h3eb75eff;
        mem[14'd6620] <= 32'h3e7799f0;
        mem[14'd6621] <= 32'h3e34b17e;
        mem[14'd6622] <= 32'h3df67077;
        mem[14'd6623] <= 32'h3e87836d;
        mem[14'd6624] <= 32'h3ea8456a;
        mem[14'd6625] <= 32'h3e03fd06;
        mem[14'd6626] <= 32'h3e595f5b;
        mem[14'd6627] <= 32'h3e9320ba;
        mem[14'd6628] <= 32'h3e8896c3;
        mem[14'd6629] <= 32'h3e81ac1c;
        mem[14'd6630] <= 32'h3eaab754;
        mem[14'd6631] <= 32'h3e317dd7;
        mem[14'd6632] <= 32'h3e4034c8;
        mem[14'd6633] <= 32'h3c3ecdc3;
        mem[14'd6634] <= 32'h3e016d92;
        mem[14'd6635] <= 32'h3d02e6f3;
        mem[14'd6636] <= 32'hbdd99a16;
        mem[14'd6637] <= 32'hbdcde41c;
        mem[14'd6638] <= 32'hbc335f8d;
        mem[14'd6639] <= 32'hbc36c7df;
        mem[14'd6640] <= 32'hbbcaab0e;
        mem[14'd6641] <= 32'h3d585750;
        mem[14'd6642] <= 32'h3dca1db0;
        mem[14'd6643] <= 32'h3e73d6f5;
        mem[14'd6644] <= 32'h3e9bb9a5;
        mem[14'd6645] <= 32'h3e5e1e5e;
        mem[14'd6646] <= 32'h3e014b59;
        mem[14'd6647] <= 32'h3db0db44;
        mem[14'd6648] <= 32'h3d87443b;
        mem[14'd6649] <= 32'h3da69b1e;
        mem[14'd6650] <= 32'hbc83a75a;
        mem[14'd6651] <= 32'h3e1bde2e;
        mem[14'd6652] <= 32'h3e96f001;
        mem[14'd6653] <= 32'h3e134bca;
        mem[14'd6654] <= 32'h3eba06f8;
        mem[14'd6655] <= 32'h3eb732bc;
        mem[14'd6656] <= 32'h3eb35b93;
        mem[14'd6657] <= 32'h3eca1571;
        mem[14'd6658] <= 32'h3e930827;
        mem[14'd6659] <= 32'h3e848113;
        mem[14'd6660] <= 32'h3e085b17;
        mem[14'd6661] <= 32'h3e4afb28;
        mem[14'd6662] <= 32'h3e161ca3;
        mem[14'd6663] <= 32'hbd229ddf;
        mem[14'd6664] <= 32'hbdb4421e;
        mem[14'd6665] <= 32'hbd63f083;
        mem[14'd6666] <= 32'hbc439cc8;
        mem[14'd6667] <= 32'h3c126fa2;
        mem[14'd6668] <= 32'h3c519a2f;
        mem[14'd6669] <= 32'h3d24f2fa;
        mem[14'd6670] <= 32'h3e0da673;
        mem[14'd6671] <= 32'h3e8f5e82;
        mem[14'd6672] <= 32'h3ea82951;
        mem[14'd6673] <= 32'h3e7ca20f;
        mem[14'd6674] <= 32'h3d80a9c8;
        mem[14'd6675] <= 32'h3d904396;
        mem[14'd6676] <= 32'hbd804214;
        mem[14'd6677] <= 32'h3d05984f;
        mem[14'd6678] <= 32'h3c567535;
        mem[14'd6679] <= 32'hbd10ca13;
        mem[14'd6680] <= 32'hbda24f20;
        mem[14'd6681] <= 32'h3e456c07;
        mem[14'd6682] <= 32'h3e9b7ab0;
        mem[14'd6683] <= 32'h3ee546f9;
        mem[14'd6684] <= 32'h3f084f8a;
        mem[14'd6685] <= 32'h3eaa080c;
        mem[14'd6686] <= 32'h3ead8d99;
        mem[14'd6687] <= 32'h3ead8232;
        mem[14'd6688] <= 32'h3ebaf16e;
        mem[14'd6689] <= 32'h3eb70c6c;
        mem[14'd6690] <= 32'h3e466380;
        mem[14'd6691] <= 32'hbde98d36;
        mem[14'd6692] <= 32'hbdf9dd0e;
        mem[14'd6693] <= 32'hbd1d20ae;
        mem[14'd6694] <= 32'h3c193644;
        mem[14'd6695] <= 32'h3b055988;
        mem[14'd6696] <= 32'hba95cfc5;
        mem[14'd6697] <= 32'h3d4de153;
        mem[14'd6698] <= 32'h3e4d1474;
        mem[14'd6699] <= 32'h3e9af01a;
        mem[14'd6700] <= 32'h3eb9bffb;
        mem[14'd6701] <= 32'h3e1fa2e5;
        mem[14'd6702] <= 32'h3c9cd00a;
        mem[14'd6703] <= 32'h3dd0d09f;
        mem[14'd6704] <= 32'h3c64521d;
        mem[14'd6705] <= 32'h3e0489a2;
        mem[14'd6706] <= 32'h3e343000;
        mem[14'd6707] <= 32'h3de65f1c;
        mem[14'd6708] <= 32'hbc986148;
        mem[14'd6709] <= 32'h3d9ca908;
        mem[14'd6710] <= 32'h3e9a05fc;
        mem[14'd6711] <= 32'h3ee4fa65;
        mem[14'd6712] <= 32'h3edd7932;
        mem[14'd6713] <= 32'h3eb7c58e;
        mem[14'd6714] <= 32'h3ee00557;
        mem[14'd6715] <= 32'h3e4f155f;
        mem[14'd6716] <= 32'h3e8c6a6c;
        mem[14'd6717] <= 32'h3e8c6b9d;
        mem[14'd6718] <= 32'h3e155521;
        mem[14'd6719] <= 32'hbdbd105d;
        mem[14'd6720] <= 32'hbddd813b;
        mem[14'd6721] <= 32'hbd45036b;
        mem[14'd6722] <= 32'hbce2cb93;
        mem[14'd6723] <= 32'h3b9bd48b;
        mem[14'd6724] <= 32'hbc12d70c;
        mem[14'd6725] <= 32'h3d4d744b;
        mem[14'd6726] <= 32'h3e4d86dc;
        mem[14'd6727] <= 32'h3eb0ec52;
        mem[14'd6728] <= 32'h3eb55613;
        mem[14'd6729] <= 32'h3e082608;
        mem[14'd6730] <= 32'h3c6be603;
        mem[14'd6731] <= 32'h3e414835;
        mem[14'd6732] <= 32'h3e845d39;
        mem[14'd6733] <= 32'hbc120a46;
        mem[14'd6734] <= 32'hbcd08eb1;
        mem[14'd6735] <= 32'hbdc44c6c;
        mem[14'd6736] <= 32'hbf066efe;
        mem[14'd6737] <= 32'hbf27f085;
        mem[14'd6738] <= 32'hbe0ce46f;
        mem[14'd6739] <= 32'h3e978777;
        mem[14'd6740] <= 32'h3ee3245f;
        mem[14'd6741] <= 32'h3ec53ae9;
        mem[14'd6742] <= 32'h3e90c57f;
        mem[14'd6743] <= 32'h3c31cdf9;
        mem[14'd6744] <= 32'h3de08cd5;
        mem[14'd6745] <= 32'h3db3f007;
        mem[14'd6746] <= 32'h3db33b56;
        mem[14'd6747] <= 32'hbd9d7a94;
        mem[14'd6748] <= 32'hbdc81d30;
        mem[14'd6749] <= 32'h3b33a73a;
        mem[14'd6750] <= 32'h3caf867f;
        mem[14'd6751] <= 32'h3c342f61;
        mem[14'd6752] <= 32'hbc87e76e;
        mem[14'd6753] <= 32'h3c263252;
        mem[14'd6754] <= 32'h3df4f15f;
        mem[14'd6755] <= 32'h3e77a6dd;
        mem[14'd6756] <= 32'h3e601cbc;
        mem[14'd6757] <= 32'h3dc9d5a3;
        mem[14'd6758] <= 32'h3dc9921e;
        mem[14'd6759] <= 32'h3d80e38a;
        mem[14'd6760] <= 32'hbcd0abe0;
        mem[14'd6761] <= 32'hbdfad120;
        mem[14'd6762] <= 32'hbd893045;
        mem[14'd6763] <= 32'hbeced646;
        mem[14'd6764] <= 32'hbf5dc79a;
        mem[14'd6765] <= 32'hbf625e93;
        mem[14'd6766] <= 32'hbe69a097;
        mem[14'd6767] <= 32'h3d926e4c;
        mem[14'd6768] <= 32'h3e5593c7;
        mem[14'd6769] <= 32'h3de4db38;
        mem[14'd6770] <= 32'h3d446390;
        mem[14'd6771] <= 32'hbcb60061;
        mem[14'd6772] <= 32'h3e2a2c22;
        mem[14'd6773] <= 32'h3d8decc3;
        mem[14'd6774] <= 32'h3cc29c61;
        mem[14'd6775] <= 32'hbd06e768;
        mem[14'd6776] <= 32'h3c248f67;
        mem[14'd6777] <= 32'h3cddf2e2;
        mem[14'd6778] <= 32'h3bfbfecb;
        mem[14'd6779] <= 32'h3b56d8d7;
        mem[14'd6780] <= 32'h3c99a50e;
        mem[14'd6781] <= 32'h3c92a475;
        mem[14'd6782] <= 32'h3d8c21b2;
        mem[14'd6783] <= 32'h3e065ed4;
        mem[14'd6784] <= 32'h3dcce12b;
        mem[14'd6785] <= 32'h3dbc69ef;
        mem[14'd6786] <= 32'hbd002560;
        mem[14'd6787] <= 32'hbd91fa72;
        mem[14'd6788] <= 32'hbdf6d307;
        mem[14'd6789] <= 32'hbe6297cd;
        mem[14'd6790] <= 32'hbe77b8ed;
        mem[14'd6791] <= 32'hbf0aa3d5;
        mem[14'd6792] <= 32'hbf5cc191;
        mem[14'd6793] <= 32'hbf1475c6;
        mem[14'd6794] <= 32'hbe2f1813;
        mem[14'd6795] <= 32'hbda1019a;
        mem[14'd6796] <= 32'h3d6ee5e9;
        mem[14'd6797] <= 32'h3e5f769d;
        mem[14'd6798] <= 32'h3eca84ae;
        mem[14'd6799] <= 32'h3ef0b441;
        mem[14'd6800] <= 32'h3e945960;
        mem[14'd6801] <= 32'h3e1343af;
        mem[14'd6802] <= 32'h3e51137b;
        mem[14'd6803] <= 32'h3e3d66be;
        mem[14'd6804] <= 32'h3c627a1c;
        mem[14'd6805] <= 32'hbc733ace;
        mem[14'd6806] <= 32'hbb83a21c;
        mem[14'd6807] <= 32'hb9178e96;
        mem[14'd6808] <= 32'hbb93e3cd;
        mem[14'd6809] <= 32'h3bbe3c17;
        mem[14'd6810] <= 32'h388d26be;
        mem[14'd6811] <= 32'h3d6784b5;
        mem[14'd6812] <= 32'h3c60a6c1;
        mem[14'd6813] <= 32'hbdb2a81b;
        mem[14'd6814] <= 32'hbd2dcfc3;
        mem[14'd6815] <= 32'hbdede972;
        mem[14'd6816] <= 32'hbe9b42dc;
        mem[14'd6817] <= 32'hbea8d8c1;
        mem[14'd6818] <= 32'hbe9a23c3;
        mem[14'd6819] <= 32'hbf065db9;
        mem[14'd6820] <= 32'hbf1a669d;
        mem[14'd6821] <= 32'hbeb75604;
        mem[14'd6822] <= 32'hbe83bef4;
        mem[14'd6823] <= 32'hbb1e8f0b;
        mem[14'd6824] <= 32'hbdb211ae;
        mem[14'd6825] <= 32'h3efe3e61;
        mem[14'd6826] <= 32'h3ef5d504;
        mem[14'd6827] <= 32'h3ebbe8f2;
        mem[14'd6828] <= 32'h3ec839ef;
        mem[14'd6829] <= 32'h3ea88ff7;
        mem[14'd6830] <= 32'h3e97a465;
        mem[14'd6831] <= 32'h3e22667e;
        mem[14'd6832] <= 32'hbc15502d;
        mem[14'd6833] <= 32'hbd4312cc;
        mem[14'd6834] <= 32'hbc16288a;
        mem[14'd6835] <= 32'hbba93afd;
        mem[14'd6836] <= 32'h3b1373b1;
        mem[14'd6837] <= 32'h3c0572dc;
        mem[14'd6838] <= 32'hba239080;
        mem[14'd6839] <= 32'hbcbcc872;
        mem[14'd6840] <= 32'h3c9f842e;
        mem[14'd6841] <= 32'hbdbb84f9;
        mem[14'd6842] <= 32'hbd52861a;
        mem[14'd6843] <= 32'h3cc818c7;
        mem[14'd6844] <= 32'hbde1f123;
        mem[14'd6845] <= 32'hbe5a45d5;
        mem[14'd6846] <= 32'hbece3895;
        mem[14'd6847] <= 32'hbf1bfffc;
        mem[14'd6848] <= 32'hbe95ff6a;
        mem[14'd6849] <= 32'hbe20ee87;
        mem[14'd6850] <= 32'hbe7a76dd;
        mem[14'd6851] <= 32'h3dc954b2;
        mem[14'd6852] <= 32'h3db939a3;
        mem[14'd6853] <= 32'h3ea12aa7;
        mem[14'd6854] <= 32'h3e36c807;
        mem[14'd6855] <= 32'h3e84ef45;
        mem[14'd6856] <= 32'h3e6d75af;
        mem[14'd6857] <= 32'h3e4e7d87;
        mem[14'd6858] <= 32'h3d5afa14;
        mem[14'd6859] <= 32'hbd2b2cbe;
        mem[14'd6860] <= 32'hbd805e28;
        mem[14'd6861] <= 32'hbd4f2522;
        mem[14'd6862] <= 32'hbac810a3;
        mem[14'd6863] <= 32'hbcba5aff;
        mem[14'd6864] <= 32'hbbbe868d;
        mem[14'd6865] <= 32'h3c747518;
        mem[14'd6866] <= 32'hbc30806a;
        mem[14'd6867] <= 32'hbcee9a24;
        mem[14'd6868] <= 32'h3ca2b4bd;
        mem[14'd6869] <= 32'hbd3ae010;
        mem[14'd6870] <= 32'hbe0fc1aa;
        mem[14'd6871] <= 32'hbe4e8bbb;
        mem[14'd6872] <= 32'hbe435a33;
        mem[14'd6873] <= 32'hbe6e493b;
        mem[14'd6874] <= 32'hbedbcd2d;
        mem[14'd6875] <= 32'hbe87e712;
        mem[14'd6876] <= 32'hbca8e0bc;
        mem[14'd6877] <= 32'h3d6d51e7;
        mem[14'd6878] <= 32'h3dd141c7;
        mem[14'd6879] <= 32'h3dc31216;
        mem[14'd6880] <= 32'hbb38a67c;
        mem[14'd6881] <= 32'hbc475055;
        mem[14'd6882] <= 32'h3d78a74a;
        mem[14'd6883] <= 32'h3d126ac7;
        mem[14'd6884] <= 32'h3db0abfb;
        mem[14'd6885] <= 32'hbc5e96c8;
        mem[14'd6886] <= 32'hbcd5f7c6;
        mem[14'd6887] <= 32'hbd754c0a;
        mem[14'd6888] <= 32'h3a9fb910;
        mem[14'd6889] <= 32'hbc1b6f0f;
        mem[14'd6890] <= 32'h3bb6a056;
        mem[14'd6891] <= 32'hbb142b27;
        mem[14'd6892] <= 32'hbbb2d1e0;
        mem[14'd6893] <= 32'h39935ac0;
        mem[14'd6894] <= 32'h3c156dfb;
        mem[14'd6895] <= 32'hbcac14c7;
        mem[14'd6896] <= 32'hbd3c3dba;
        mem[14'd6897] <= 32'hbe056f36;
        mem[14'd6898] <= 32'hbeaa6ebb;
        mem[14'd6899] <= 32'hbea38e05;
        mem[14'd6900] <= 32'hbe9e7585;
        mem[14'd6901] <= 32'hbeae4ce1;
        mem[14'd6902] <= 32'hbeb6faa1;
        mem[14'd6903] <= 32'hbe32d50c;
        mem[14'd6904] <= 32'hbdd04deb;
        mem[14'd6905] <= 32'h3d7819d1;
        mem[14'd6906] <= 32'h3cfadcca;
        mem[14'd6907] <= 32'hbd54a230;
        mem[14'd6908] <= 32'hbe3f9ab7;
        mem[14'd6909] <= 32'hbdcf57d3;
        mem[14'd6910] <= 32'hbd92d392;
        mem[14'd6911] <= 32'hbd730d71;
        mem[14'd6912] <= 32'hbd9433a3;
        mem[14'd6913] <= 32'hbe237dde;
        mem[14'd6914] <= 32'hbe3c653d;
        mem[14'd6915] <= 32'hbe3bb3e9;
        mem[14'd6916] <= 32'hbdad5d17;
        mem[14'd6917] <= 32'hbc56aff3;
        mem[14'd6918] <= 32'h3cf69797;
        mem[14'd6919] <= 32'hba431cac;
        mem[14'd6920] <= 32'hbcbad705;
        mem[14'd6921] <= 32'h3c8d8090;
        mem[14'd6922] <= 32'h3c30c16c;
        mem[14'd6923] <= 32'hbd602924;
        mem[14'd6924] <= 32'hbdcb8ecb;
        mem[14'd6925] <= 32'hbe51a34e;
        mem[14'd6926] <= 32'hbeaaf5aa;
        mem[14'd6927] <= 32'hbec87ada;
        mem[14'd6928] <= 32'hbea7c7cb;
        mem[14'd6929] <= 32'hbe95f729;
        mem[14'd6930] <= 32'hbeb2143b;
        mem[14'd6931] <= 32'hbe55a790;
        mem[14'd6932] <= 32'hbdac534e;
        mem[14'd6933] <= 32'hbd28c779;
        mem[14'd6934] <= 32'h3db40403;
        mem[14'd6935] <= 32'hbe0e6fa9;
        mem[14'd6936] <= 32'hbe868f6e;
        mem[14'd6937] <= 32'hbe84b37c;
        mem[14'd6938] <= 32'hbe9c23d0;
        mem[14'd6939] <= 32'hbe45cd46;
        mem[14'd6940] <= 32'hbe950493;
        mem[14'd6941] <= 32'hbebcb7f9;
        mem[14'd6942] <= 32'hbeac9c01;
        mem[14'd6943] <= 32'hbe6ece8e;
        mem[14'd6944] <= 32'hbd85249a;
        mem[14'd6945] <= 32'hbcd3a0a0;
        mem[14'd6946] <= 32'hbc1a16ba;
        mem[14'd6947] <= 32'hbbcde2a4;
        mem[14'd6948] <= 32'h3c246802;
        mem[14'd6949] <= 32'hbbd6b68c;
        mem[14'd6950] <= 32'hbc201707;
        mem[14'd6951] <= 32'hbd45285a;
        mem[14'd6952] <= 32'hbe185c4c;
        mem[14'd6953] <= 32'hbe75cda8;
        mem[14'd6954] <= 32'hbeb963e5;
        mem[14'd6955] <= 32'hbecaed0f;
        mem[14'd6956] <= 32'hbe991b7d;
        mem[14'd6957] <= 32'hbe932d21;
        mem[14'd6958] <= 32'hbe8e1545;
        mem[14'd6959] <= 32'hbe6985bd;
        mem[14'd6960] <= 32'hbd387632;
        mem[14'd6961] <= 32'h3bd4d184;
        mem[14'd6962] <= 32'h3d13ca62;
        mem[14'd6963] <= 32'hbe22492e;
        mem[14'd6964] <= 32'hbe9a136e;
        mem[14'd6965] <= 32'hbeaa378d;
        mem[14'd6966] <= 32'hbef9703c;
        mem[14'd6967] <= 32'hbeb7dc06;
        mem[14'd6968] <= 32'hbee43141;
        mem[14'd6969] <= 32'hbee7d457;
        mem[14'd6970] <= 32'hbec7f452;
        mem[14'd6971] <= 32'hbe3d1317;
        mem[14'd6972] <= 32'hbd3f1ded;
        mem[14'd6973] <= 32'hbcd5aaf3;
        mem[14'd6974] <= 32'h3c9b8623;
        mem[14'd6975] <= 32'hbcb509a7;
        mem[14'd6976] <= 32'h3b9b7f63;
        mem[14'd6977] <= 32'h3b123a0a;
        mem[14'd6978] <= 32'hbd121239;
        mem[14'd6979] <= 32'hbdb2f09a;
        mem[14'd6980] <= 32'hbe24cec4;
        mem[14'd6981] <= 32'hbe575c6f;
        mem[14'd6982] <= 32'hbe9e7dd6;
        mem[14'd6983] <= 32'hbea3e434;
        mem[14'd6984] <= 32'hbe5d25b3;
        mem[14'd6985] <= 32'hbe867f9a;
        mem[14'd6986] <= 32'hbe5a8888;
        mem[14'd6987] <= 32'hbe2c22f0;
        mem[14'd6988] <= 32'hbdb274aa;
        mem[14'd6989] <= 32'hbe02545e;
        mem[14'd6990] <= 32'hbe1dffa4;
        mem[14'd6991] <= 32'hbe03d955;
        mem[14'd6992] <= 32'hbe0b82d1;
        mem[14'd6993] <= 32'hbe91b173;
        mem[14'd6994] <= 32'hbebb38cc;
        mem[14'd6995] <= 32'hbecbf2d8;
        mem[14'd6996] <= 32'hbed81607;
        mem[14'd6997] <= 32'hbec3bd23;
        mem[14'd6998] <= 32'hbea6d0c6;
        mem[14'd6999] <= 32'hbe4c7ba4;
        mem[14'd7000] <= 32'hbd107f2b;
        mem[14'd7001] <= 32'hbc17f326;
        mem[14'd7002] <= 32'h3c1d7e5f;
        mem[14'd7003] <= 32'h3c539f0f;
        mem[14'd7004] <= 32'h3c2ad638;
        mem[14'd7005] <= 32'h3a00a18e;
        mem[14'd7006] <= 32'hbceffd6f;
        mem[14'd7007] <= 32'hbd9061a7;
        mem[14'd7008] <= 32'hbdb88798;
        mem[14'd7009] <= 32'hbd4aa26e;
        mem[14'd7010] <= 32'hbd8f19a7;
        mem[14'd7011] <= 32'hbbbc1756;
        mem[14'd7012] <= 32'hbd97b20b;
        mem[14'd7013] <= 32'hbe21699f;
        mem[14'd7014] <= 32'hbe0a02f5;
        mem[14'd7015] <= 32'hbe555aac;
        mem[14'd7016] <= 32'hbdbd2ac9;
        mem[14'd7017] <= 32'hbe81b9be;
        mem[14'd7018] <= 32'hbdf5f1fd;
        mem[14'd7019] <= 32'hbd28ab96;
        mem[14'd7020] <= 32'hbd7be0da;
        mem[14'd7021] <= 32'hbe7b2425;
        mem[14'd7022] <= 32'hbe920907;
        mem[14'd7023] <= 32'hbe974f52;
        mem[14'd7024] <= 32'hbebc10c7;
        mem[14'd7025] <= 32'hbeaf7844;
        mem[14'd7026] <= 32'hbe919882;
        mem[14'd7027] <= 32'hbe382b0a;
        mem[14'd7028] <= 32'hbcb620c7;
        mem[14'd7029] <= 32'hbb923f44;
        mem[14'd7030] <= 32'h3b7995b0;
        mem[14'd7031] <= 32'h3c0c31f9;
        mem[14'd7032] <= 32'h3c4538bd;
        mem[14'd7033] <= 32'hbc3303aa;
        mem[14'd7034] <= 32'hbce42e74;
        mem[14'd7035] <= 32'hbd23396c;
        mem[14'd7036] <= 32'hba258b59;
        mem[14'd7037] <= 32'h3dcc3efb;
        mem[14'd7038] <= 32'h3e4f35f9;
        mem[14'd7039] <= 32'h3e77c9b9;
        mem[14'd7040] <= 32'hbdccbc15;
        mem[14'd7041] <= 32'hbdb698d8;
        mem[14'd7042] <= 32'hbdd29b26;
        mem[14'd7043] <= 32'hbe483b4a;
        mem[14'd7044] <= 32'hbe52e1e9;
        mem[14'd7045] <= 32'hbe46dd3b;
        mem[14'd7046] <= 32'hbd97af7e;
        mem[14'd7047] <= 32'h3c5c59c9;
        mem[14'd7048] <= 32'hbdbfed29;
        mem[14'd7049] <= 32'hbdf534de;
        mem[14'd7050] <= 32'hbe66603d;
        mem[14'd7051] <= 32'hbe9b6b90;
        mem[14'd7052] <= 32'hbeac3c67;
        mem[14'd7053] <= 32'hbea14304;
        mem[14'd7054] <= 32'hbe5d6411;
        mem[14'd7055] <= 32'hbe36915c;
        mem[14'd7056] <= 32'hbd50d603;
        mem[14'd7057] <= 32'h3b8d6214;
        mem[14'd7058] <= 32'hbb07a998;
        mem[14'd7059] <= 32'hbb91f0c6;
        mem[14'd7060] <= 32'hbb7e6ecf;
        mem[14'd7061] <= 32'h3b107f88;
        mem[14'd7062] <= 32'h3c4a1525;
        mem[14'd7063] <= 32'h3b983544;
        mem[14'd7064] <= 32'h3daa1193;
        mem[14'd7065] <= 32'h3e839bcf;
        mem[14'd7066] <= 32'h3e9d1dde;
        mem[14'd7067] <= 32'h3e895e83;
        mem[14'd7068] <= 32'h3e285c65;
        mem[14'd7069] <= 32'h3da468a3;
        mem[14'd7070] <= 32'h3de8bba4;
        mem[14'd7071] <= 32'h3d97ac77;
        mem[14'd7072] <= 32'h3d693ad4;
        mem[14'd7073] <= 32'h3ddb853e;
        mem[14'd7074] <= 32'h3d7a3596;
        mem[14'd7075] <= 32'h3d80bb54;
        mem[14'd7076] <= 32'hbc1b959a;
        mem[14'd7077] <= 32'h3c791551;
        mem[14'd7078] <= 32'hbdf8eb6f;
        mem[14'd7079] <= 32'hbe186569;
        mem[14'd7080] <= 32'hbe34b454;
        mem[14'd7081] <= 32'hbe3bc0f6;
        mem[14'd7082] <= 32'hbe195dea;
        mem[14'd7083] <= 32'hbe0d5f2b;
        mem[14'd7084] <= 32'hbd83e9ab;
        mem[14'd7085] <= 32'hbbea48ad;
        mem[14'd7086] <= 32'hbb572245;
        mem[14'd7087] <= 32'h3cc129e9;
        mem[14'd7088] <= 32'hbae5ed06;
        mem[14'd7089] <= 32'h3c2c273d;
        mem[14'd7090] <= 32'h3ba83e96;
        mem[14'd7091] <= 32'h3bf9a73e;
        mem[14'd7092] <= 32'h3d9c2a40;
        mem[14'd7093] <= 32'h3dc3a33e;
        mem[14'd7094] <= 32'h3ddc9dd9;
        mem[14'd7095] <= 32'h3e37dc87;
        mem[14'd7096] <= 32'h3e964385;
        mem[14'd7097] <= 32'h3ea57b25;
        mem[14'd7098] <= 32'h3e80c4ba;
        mem[14'd7099] <= 32'h3ec22c1b;
        mem[14'd7100] <= 32'h3ea2ea13;
        mem[14'd7101] <= 32'h3e77b9a9;
        mem[14'd7102] <= 32'h3e803179;
        mem[14'd7103] <= 32'h3e6baf4b;
        mem[14'd7104] <= 32'h3e4a958d;
        mem[14'd7105] <= 32'h3e4cfd17;
        mem[14'd7106] <= 32'h3e1ec57b;
        mem[14'd7107] <= 32'h3d2caa97;
        mem[14'd7108] <= 32'hbdabf035;
        mem[14'd7109] <= 32'hbd88d13f;
        mem[14'd7110] <= 32'hbd106089;
        mem[14'd7111] <= 32'hbcfed4b1;
        mem[14'd7112] <= 32'hbb72bd5d;
        mem[14'd7113] <= 32'h39c46102;
        mem[14'd7114] <= 32'hb91b1c0c;
        mem[14'd7115] <= 32'h3a791a22;
        mem[14'd7116] <= 32'hbb0cacf7;
        mem[14'd7117] <= 32'hbaebabbc;
        mem[14'd7118] <= 32'h3c869886;
        mem[14'd7119] <= 32'hbce32661;
        mem[14'd7120] <= 32'hbccc34a9;
        mem[14'd7121] <= 32'hbd03fae5;
        mem[14'd7122] <= 32'hbd67c61a;
        mem[14'd7123] <= 32'hbb0a9b0c;
        mem[14'd7124] <= 32'h3d993d4d;
        mem[14'd7125] <= 32'h3ddbeaf5;
        mem[14'd7126] <= 32'h3e131e8f;
        mem[14'd7127] <= 32'h3de1ec56;
        mem[14'd7128] <= 32'h3dc74e6f;
        mem[14'd7129] <= 32'h3e630a39;
        mem[14'd7130] <= 32'h3e85d6a6;
        mem[14'd7131] <= 32'h3e9512d8;
        mem[14'd7132] <= 32'h3e673dac;
        mem[14'd7133] <= 32'h3e70b1dd;
        mem[14'd7134] <= 32'h3e65c8ea;
        mem[14'd7135] <= 32'h3e08b6f4;
        mem[14'd7136] <= 32'h3c02de4f;
        mem[14'd7137] <= 32'h3cf4f3a7;
        mem[14'd7138] <= 32'h3c4eb2af;
        mem[14'd7139] <= 32'h3ba53d0f;
        mem[14'd7140] <= 32'h3b4e6462;
        mem[14'd7141] <= 32'hba92acf6;
        mem[14'd7142] <= 32'h3a96b37a;
        mem[14'd7143] <= 32'h3acfdfb8;
        mem[14'd7144] <= 32'hbbb54b21;
        mem[14'd7145] <= 32'hbc0106f6;
        mem[14'd7146] <= 32'hbc4c6b1c;
        mem[14'd7147] <= 32'h3c757beb;
        mem[14'd7148] <= 32'h3bb3b33d;
        mem[14'd7149] <= 32'h3c540977;
        mem[14'd7150] <= 32'hbcaf9a43;
        mem[14'd7151] <= 32'h3c43e9e4;
        mem[14'd7152] <= 32'h3c398e2b;
        mem[14'd7153] <= 32'h3c90e0e8;
        mem[14'd7154] <= 32'h3cfd31f9;
        mem[14'd7155] <= 32'h3cf00841;
        mem[14'd7156] <= 32'h3c88b3ec;
        mem[14'd7157] <= 32'h3db5fdbe;
        mem[14'd7158] <= 32'h3db9cb2a;
        mem[14'd7159] <= 32'h3d9043e9;
        mem[14'd7160] <= 32'h3d83a4ef;
        mem[14'd7161] <= 32'h3dc3b7c1;
        mem[14'd7162] <= 32'h3da3bd12;
        mem[14'd7163] <= 32'h3d7a0a84;
        mem[14'd7164] <= 32'h3cc1b4f2;
        mem[14'd7165] <= 32'h3d097f3c;
        mem[14'd7166] <= 32'h3c968562;
        mem[14'd7167] <= 32'h3b16410c;
        mem[14'd7168] <= 32'hbb81f103;
        mem[14'd7169] <= 32'h38ab21a2;
        mem[14'd7170] <= 32'h3ca69904;
        mem[14'd7171] <= 32'h3c0dffd9;
        mem[14'd7172] <= 32'hbc460a5c;
        mem[14'd7173] <= 32'hbccb66c2;
        mem[14'd7174] <= 32'h3b931ac9;
        mem[14'd7175] <= 32'hbc3a6ae6;
        mem[14'd7176] <= 32'hbba93713;
        mem[14'd7177] <= 32'hbc24dbe2;
        mem[14'd7178] <= 32'h39c2fc6b;
        mem[14'd7179] <= 32'h3ba2e236;
        mem[14'd7180] <= 32'hbb08c891;
        mem[14'd7181] <= 32'h3c4944be;
        mem[14'd7182] <= 32'h3c723fd9;
        mem[14'd7183] <= 32'hbbdeca9d;
        mem[14'd7184] <= 32'hbb42d969;
        mem[14'd7185] <= 32'h3c06f7b6;
        mem[14'd7186] <= 32'hbb88cad1;
        mem[14'd7187] <= 32'h3bebde1e;
        mem[14'd7188] <= 32'hbba66a77;
        mem[14'd7189] <= 32'hbce470fc;
        mem[14'd7190] <= 32'h3c70d23d;
        mem[14'd7191] <= 32'h3bd2ad09;
        mem[14'd7192] <= 32'h3a6c1f39;
        mem[14'd7193] <= 32'h3c34d241;
        mem[14'd7194] <= 32'h3c94e8c7;
        mem[14'd7195] <= 32'h3c62a7b0;
        mem[14'd7196] <= 32'hbc07cf35;
        mem[14'd7197] <= 32'h3c181572;
        mem[14'd7198] <= 32'hbcaf632a;
        mem[14'd7199] <= 32'hbb292573;
        mem[14'd7200] <= 32'hbbf7b7d9;
        mem[14'd7201] <= 32'hbc23acb7;
        mem[14'd7202] <= 32'h3b10ec73;
        mem[14'd7203] <= 32'hbbc1c224;
        mem[14'd7204] <= 32'hbbda9177;
        mem[14'd7205] <= 32'hbba7fe22;
        mem[14'd7206] <= 32'hbc780d60;
        mem[14'd7207] <= 32'h3bb9dccf;
        mem[14'd7208] <= 32'h3beb6fd5;
        mem[14'd7209] <= 32'h3c45a6df;
        mem[14'd7210] <= 32'h3c26519a;
        mem[14'd7211] <= 32'hbbb4f503;
        mem[14'd7212] <= 32'h39879d89;
        mem[14'd7213] <= 32'h3aab53e3;
        mem[14'd7214] <= 32'hbc244c38;
        mem[14'd7215] <= 32'hbc0ceb0c;
        mem[14'd7216] <= 32'h3c4f3f06;
        mem[14'd7217] <= 32'hbb34e726;
        mem[14'd7218] <= 32'hba020033;
        mem[14'd7219] <= 32'hba1dd3a0;
        mem[14'd7220] <= 32'hbacb823f;
        mem[14'd7221] <= 32'h3bb64fcd;
        mem[14'd7222] <= 32'hbbc382aa;
        mem[14'd7223] <= 32'hbc5ad549;
        mem[14'd7224] <= 32'h3c563720;
        mem[14'd7225] <= 32'hbc11fb00;
        mem[14'd7226] <= 32'h3bf449f2;
        mem[14'd7227] <= 32'h3b38ab00;
        mem[14'd7228] <= 32'hbc6bb8dc;
        mem[14'd7229] <= 32'hbac0281e;
        mem[14'd7230] <= 32'hbabd9912;
        mem[14'd7231] <= 32'hbb83e3ca;
        mem[14'd7232] <= 32'h3bbd1363;
        mem[14'd7233] <= 32'h3bd2428c;
        mem[14'd7234] <= 32'hbbf75cd8;
        mem[14'd7235] <= 32'hbc49a651;
        mem[14'd7236] <= 32'hbc241b81;
        mem[14'd7237] <= 32'hbbf94599;
        mem[14'd7238] <= 32'hbc83479d;
        mem[14'd7239] <= 32'hbc5216bd;
        mem[14'd7240] <= 32'hbc9952f2;
        mem[14'd7241] <= 32'hbcc73da5;
        mem[14'd7242] <= 32'hbd2c2070;
        mem[14'd7243] <= 32'hbd962d4b;
        mem[14'd7244] <= 32'hbd4c24ec;
        mem[14'd7245] <= 32'hbd16a4a4;
        mem[14'd7246] <= 32'hbc646224;
        mem[14'd7247] <= 32'hbcc8d2ae;
        mem[14'd7248] <= 32'h3ba4d1ed;
        mem[14'd7249] <= 32'hbbd3faad;
        mem[14'd7250] <= 32'hbc26cf7d;
        mem[14'd7251] <= 32'hbbc84de5;
        mem[14'd7252] <= 32'hbc97ee9a;
        mem[14'd7253] <= 32'h3b1a1c83;
        mem[14'd7254] <= 32'h3b89df9f;
        mem[14'd7255] <= 32'h3b7c5880;
        mem[14'd7256] <= 32'h3c2d433b;
        mem[14'd7257] <= 32'h3c4fa54a;
        mem[14'd7258] <= 32'h3c09a42f;
        mem[14'd7259] <= 32'h3c6ba699;
        mem[14'd7260] <= 32'hbc9d0626;
        mem[14'd7261] <= 32'hba91ac41;
        mem[14'd7262] <= 32'h3b9fd162;
        mem[14'd7263] <= 32'hbb897c93;
        mem[14'd7264] <= 32'hbcd2178b;
        mem[14'd7265] <= 32'hbd1c68c6;
        mem[14'd7266] <= 32'hbd00aaa3;
        mem[14'd7267] <= 32'hbd9e7df5;
        mem[14'd7268] <= 32'hbd971026;
        mem[14'd7269] <= 32'hbdabe720;
        mem[14'd7270] <= 32'hbdda0746;
        mem[14'd7271] <= 32'hbdf2463c;
        mem[14'd7272] <= 32'hbdcf6724;
        mem[14'd7273] <= 32'hbd9aa245;
        mem[14'd7274] <= 32'hbc6c5de7;
        mem[14'd7275] <= 32'hbda3fe4b;
        mem[14'd7276] <= 32'hbd147f7c;
        mem[14'd7277] <= 32'h3c000f10;
        mem[14'd7278] <= 32'h3cbd00b8;
        mem[14'd7279] <= 32'h3cb77340;
        mem[14'd7280] <= 32'h3c30de6f;
        mem[14'd7281] <= 32'h3bfbf1bb;
        mem[14'd7282] <= 32'hbc49d0ce;
        mem[14'd7283] <= 32'h3bc4ad78;
        mem[14'd7284] <= 32'hbbf005bb;
        mem[14'd7285] <= 32'h3bdb01ab;
        mem[14'd7286] <= 32'hbbc094a3;
        mem[14'd7287] <= 32'hbc7e04a4;
        mem[14'd7288] <= 32'hbb32ece3;
        mem[14'd7289] <= 32'hbc080b98;
        mem[14'd7290] <= 32'hbd100e9e;
        mem[14'd7291] <= 32'hbd0d66de;
        mem[14'd7292] <= 32'h3ca2f5a0;
        mem[14'd7293] <= 32'h3d42ca43;
        mem[14'd7294] <= 32'h3d3ff183;
        mem[14'd7295] <= 32'h3dea4011;
        mem[14'd7296] <= 32'h3e586f5f;
        mem[14'd7297] <= 32'h3e22cc6f;
        mem[14'd7298] <= 32'h3e933fd1;
        mem[14'd7299] <= 32'h3e81ba76;
        mem[14'd7300] <= 32'h3e6c19fd;
        mem[14'd7301] <= 32'h3dc80064;
        mem[14'd7302] <= 32'h3d838634;
        mem[14'd7303] <= 32'h3d107382;
        mem[14'd7304] <= 32'h3da067d0;
        mem[14'd7305] <= 32'hbc9b9c73;
        mem[14'd7306] <= 32'hbd51d98f;
        mem[14'd7307] <= 32'hbd781a67;
        mem[14'd7308] <= 32'h3cd2835c;
        mem[14'd7309] <= 32'h3d1ff83d;
        mem[14'd7310] <= 32'h3cebfaa9;
        mem[14'd7311] <= 32'h3c8167d7;
        mem[14'd7312] <= 32'h3c7f9080;
        mem[14'd7313] <= 32'h3bd254be;
        mem[14'd7314] <= 32'hbbd956e1;
        mem[14'd7315] <= 32'h3b0b91f1;
        mem[14'd7316] <= 32'hbd1e29d3;
        mem[14'd7317] <= 32'hbd437e3f;
        mem[14'd7318] <= 32'hbd87de9b;
        mem[14'd7319] <= 32'hbd2741a5;
        mem[14'd7320] <= 32'hbd1ade33;
        mem[14'd7321] <= 32'h3d1e2227;
        mem[14'd7322] <= 32'hbd64ba9b;
        mem[14'd7323] <= 32'h3e134fbf;
        mem[14'd7324] <= 32'h3e7b2c35;
        mem[14'd7325] <= 32'h3e1f5ff1;
        mem[14'd7326] <= 32'h3e3753ef;
        mem[14'd7327] <= 32'h3def2c35;
        mem[14'd7328] <= 32'h3e304ece;
        mem[14'd7329] <= 32'h3e7a38b7;
        mem[14'd7330] <= 32'hbc82f24c;
        mem[14'd7331] <= 32'h3dcff98f;
        mem[14'd7332] <= 32'h3e2370dd;
        mem[14'd7333] <= 32'h3d2b9831;
        mem[14'd7334] <= 32'hbd9af074;
        mem[14'd7335] <= 32'hbe091666;
        mem[14'd7336] <= 32'hbc81c72b;
        mem[14'd7337] <= 32'h3d925f9e;
        mem[14'd7338] <= 32'h3bdb076f;
        mem[14'd7339] <= 32'h3c01e9f0;
        mem[14'd7340] <= 32'hbc2373e5;
        mem[14'd7341] <= 32'h3a45ddb6;
        mem[14'd7342] <= 32'hbc475b0b;
        mem[14'd7343] <= 32'hbcce981e;
        mem[14'd7344] <= 32'hbd63ca0c;
        mem[14'd7345] <= 32'hbd9d3d96;
        mem[14'd7346] <= 32'hbdecc0dd;
        mem[14'd7347] <= 32'hbd731754;
        mem[14'd7348] <= 32'h3c90e00a;
        mem[14'd7349] <= 32'h3c087833;
        mem[14'd7350] <= 32'hbd5b8521;
        mem[14'd7351] <= 32'h3cbe955b;
        mem[14'd7352] <= 32'h3e3bbed9;
        mem[14'd7353] <= 32'h3db35751;
        mem[14'd7354] <= 32'h3d37b8fe;
        mem[14'd7355] <= 32'h3e8a449a;
        mem[14'd7356] <= 32'h3dcd221d;
        mem[14'd7357] <= 32'h3df4cdda;
        mem[14'd7358] <= 32'hbdc6317c;
        mem[14'd7359] <= 32'h3e3962d1;
        mem[14'd7360] <= 32'h3dd0d83b;
        mem[14'd7361] <= 32'h3bac6d9f;
        mem[14'd7362] <= 32'hbc42fca2;
        mem[14'd7363] <= 32'h3e0e0451;
        mem[14'd7364] <= 32'h3d77c9ac;
        mem[14'd7365] <= 32'h3dc2b394;
        mem[14'd7366] <= 32'hbb29c040;
        mem[14'd7367] <= 32'hbc052e76;
        mem[14'd7368] <= 32'h3a680fd5;
        mem[14'd7369] <= 32'hbc0a28c4;
        mem[14'd7370] <= 32'h3c0413f6;
        mem[14'd7371] <= 32'hbc2a2c27;
        mem[14'd7372] <= 32'hbd2cfedc;
        mem[14'd7373] <= 32'hbd0fd906;
        mem[14'd7374] <= 32'hbd650d03;
        mem[14'd7375] <= 32'h3d103329;
        mem[14'd7376] <= 32'h3e01b312;
        mem[14'd7377] <= 32'h3c1965ec;
        mem[14'd7378] <= 32'h3cbc6c71;
        mem[14'd7379] <= 32'hbdc455f2;
        mem[14'd7380] <= 32'hbd94d8d8;
        mem[14'd7381] <= 32'hbd5459b5;
        mem[14'd7382] <= 32'hbe64d8dd;
        mem[14'd7383] <= 32'h3e21dae0;
        mem[14'd7384] <= 32'h3d22f430;
        mem[14'd7385] <= 32'hbe07bdfc;
        mem[14'd7386] <= 32'h3d799a48;
        mem[14'd7387] <= 32'h3b80d8e5;
        mem[14'd7388] <= 32'hbc9bb579;
        mem[14'd7389] <= 32'h3de99e3a;
        mem[14'd7390] <= 32'h3d25fa2a;
        mem[14'd7391] <= 32'h3e90e0b9;
        mem[14'd7392] <= 32'h3e87e1bc;
        mem[14'd7393] <= 32'h3d4f5147;
        mem[14'd7394] <= 32'h3b8706c5;
        mem[14'd7395] <= 32'hbc0e2703;
        mem[14'd7396] <= 32'hbc2aa928;
        mem[14'd7397] <= 32'h3acf60cc;
        mem[14'd7398] <= 32'hbc3a68ee;
        mem[14'd7399] <= 32'hbc6c4734;
        mem[14'd7400] <= 32'hbbb5e2dc;
        mem[14'd7401] <= 32'h3cb97389;
        mem[14'd7402] <= 32'h3e0698ef;
        mem[14'd7403] <= 32'h3e2fcf2d;
        mem[14'd7404] <= 32'h3d934377;
        mem[14'd7405] <= 32'h3e243ed3;
        mem[14'd7406] <= 32'h3da30706;
        mem[14'd7407] <= 32'hbab94b2d;
        mem[14'd7408] <= 32'h3e3d3dac;
        mem[14'd7409] <= 32'h3e3c03a9;
        mem[14'd7410] <= 32'hbe111684;
        mem[14'd7411] <= 32'hbdb57c34;
        mem[14'd7412] <= 32'h3dfb5eb9;
        mem[14'd7413] <= 32'hbd81e56b;
        mem[14'd7414] <= 32'h3da87613;
        mem[14'd7415] <= 32'h3dff1007;
        mem[14'd7416] <= 32'h3d327b4b;
        mem[14'd7417] <= 32'h3db4c13a;
        mem[14'd7418] <= 32'h3e1b89a4;
        mem[14'd7419] <= 32'h3ea5fa57;
        mem[14'd7420] <= 32'h3ec2063d;
        mem[14'd7421] <= 32'h3dd1e263;
        mem[14'd7422] <= 32'h3db09cb9;
        mem[14'd7423] <= 32'h3cd59cd4;
        mem[14'd7424] <= 32'h3b64793b;
        mem[14'd7425] <= 32'h3c7279fb;
        mem[14'd7426] <= 32'hbc8b5ba5;
        mem[14'd7427] <= 32'hbcd8bb0a;
        mem[14'd7428] <= 32'hbc1fe5ae;
        mem[14'd7429] <= 32'h3da7490b;
        mem[14'd7430] <= 32'h3e32a247;
        mem[14'd7431] <= 32'h3dfcbdbc;
        mem[14'd7432] <= 32'h3e177087;
        mem[14'd7433] <= 32'h3e441698;
        mem[14'd7434] <= 32'h3e05aa04;
        mem[14'd7435] <= 32'h3e026efb;
        mem[14'd7436] <= 32'h3ce78114;
        mem[14'd7437] <= 32'h3c8a5d60;
        mem[14'd7438] <= 32'hbe496f2f;
        mem[14'd7439] <= 32'hbed145da;
        mem[14'd7440] <= 32'hbe19abc5;
        mem[14'd7441] <= 32'h3ca32392;
        mem[14'd7442] <= 32'hbd310000;
        mem[14'd7443] <= 32'h3df48c79;
        mem[14'd7444] <= 32'h3dcacb21;
        mem[14'd7445] <= 32'h3e1aacac;
        mem[14'd7446] <= 32'h3e5f4e24;
        mem[14'd7447] <= 32'h3ea2cedd;
        mem[14'd7448] <= 32'h3e44968d;
        mem[14'd7449] <= 32'h3d0c568d;
        mem[14'd7450] <= 32'h3d5e22d4;
        mem[14'd7451] <= 32'hbcc642e1;
        mem[14'd7452] <= 32'hbba82e39;
        mem[14'd7453] <= 32'h3af8aca7;
        mem[14'd7454] <= 32'hbb9982d2;
        mem[14'd7455] <= 32'hbd6141e6;
        mem[14'd7456] <= 32'h3dc3b51e;
        mem[14'd7457] <= 32'h3de206fa;
        mem[14'd7458] <= 32'h3e2b30a4;
        mem[14'd7459] <= 32'h3e3c2b5b;
        mem[14'd7460] <= 32'h3e146e01;
        mem[14'd7461] <= 32'h3e82285f;
        mem[14'd7462] <= 32'h3ea24397;
        mem[14'd7463] <= 32'h3e506fc0;
        mem[14'd7464] <= 32'h3e4ea369;
        mem[14'd7465] <= 32'h3cea11fe;
        mem[14'd7466] <= 32'hbcaad63b;
        mem[14'd7467] <= 32'hbe9be9b4;
        mem[14'd7468] <= 32'hbe8d957b;
        mem[14'd7469] <= 32'hbe2e9548;
        mem[14'd7470] <= 32'h3daa9cac;
        mem[14'd7471] <= 32'h3e4b8dc6;
        mem[14'd7472] <= 32'h3debeb03;
        mem[14'd7473] <= 32'h3e1ebb39;
        mem[14'd7474] <= 32'h3e4653d4;
        mem[14'd7475] <= 32'h3e83b4ae;
        mem[14'd7476] <= 32'hbb9efd1a;
        mem[14'd7477] <= 32'hbdb6ac6d;
        mem[14'd7478] <= 32'h3cb18923;
        mem[14'd7479] <= 32'h3ab41c3e;
        mem[14'd7480] <= 32'h3b164719;
        mem[14'd7481] <= 32'hbcaf3f9d;
        mem[14'd7482] <= 32'hbb29b39a;
        mem[14'd7483] <= 32'hbccab09a;
        mem[14'd7484] <= 32'h3dad8f03;
        mem[14'd7485] <= 32'h3e42c445;
        mem[14'd7486] <= 32'h3e38083d;
        mem[14'd7487] <= 32'h3eb1eb67;
        mem[14'd7488] <= 32'h3e8826f7;
        mem[14'd7489] <= 32'h3e9c472a;
        mem[14'd7490] <= 32'h3e63103b;
        mem[14'd7491] <= 32'h3e1180ac;
        mem[14'd7492] <= 32'h3e47a181;
        mem[14'd7493] <= 32'h3eb1fb81;
        mem[14'd7494] <= 32'h3ededc75;
        mem[14'd7495] <= 32'hbbf2f00b;
        mem[14'd7496] <= 32'hbe3e3e6d;
        mem[14'd7497] <= 32'hbe36616f;
        mem[14'd7498] <= 32'hbde470d8;
        mem[14'd7499] <= 32'h3c993526;
        mem[14'd7500] <= 32'h3d1fb8f4;
        mem[14'd7501] <= 32'h3dc7df7e;
        mem[14'd7502] <= 32'h3e9bf603;
        mem[14'd7503] <= 32'h3eb20171;
        mem[14'd7504] <= 32'h3e82eada;
        mem[14'd7505] <= 32'h3cb47c79;
        mem[14'd7506] <= 32'h3db757a7;
        mem[14'd7507] <= 32'h3c316e7d;
        mem[14'd7508] <= 32'hb8427af0;
        mem[14'd7509] <= 32'hbc870563;
        mem[14'd7510] <= 32'hbc638c2a;
        mem[14'd7511] <= 32'h3d0a7a48;
        mem[14'd7512] <= 32'h3d8d8218;
        mem[14'd7513] <= 32'h3e5ecafe;
        mem[14'd7514] <= 32'h3df4e0e7;
        mem[14'd7515] <= 32'h3e20467d;
        mem[14'd7516] <= 32'h3cd3376d;
        mem[14'd7517] <= 32'h3e0c7d19;
        mem[14'd7518] <= 32'hbdc4b4fb;
        mem[14'd7519] <= 32'hbd149169;
        mem[14'd7520] <= 32'h3de7403d;
        mem[14'd7521] <= 32'h3ecb9b40;
        mem[14'd7522] <= 32'h3e88c59f;
        mem[14'd7523] <= 32'h3d8b787f;
        mem[14'd7524] <= 32'h3c8fa1ef;
        mem[14'd7525] <= 32'hbbcb4344;
        mem[14'd7526] <= 32'hbd6aef89;
        mem[14'd7527] <= 32'h3e12686b;
        mem[14'd7528] <= 32'h3e3ba4ff;
        mem[14'd7529] <= 32'h3ea6297b;
        mem[14'd7530] <= 32'h3eb3b090;
        mem[14'd7531] <= 32'h3ed8d6aa;
        mem[14'd7532] <= 32'h3e99fe69;
        mem[14'd7533] <= 32'h3d803cc7;
        mem[14'd7534] <= 32'h3d16021f;
        mem[14'd7535] <= 32'hbbf9812e;
        mem[14'd7536] <= 32'h3c6030aa;
        mem[14'd7537] <= 32'hbb89b37c;
        mem[14'd7538] <= 32'hbc1d44d7;
        mem[14'd7539] <= 32'hbbad2ca1;
        mem[14'd7540] <= 32'hbc78bf6b;
        mem[14'd7541] <= 32'h3d4635f7;
        mem[14'd7542] <= 32'hbc2b0705;
        mem[14'd7543] <= 32'h3ba0eeaf;
        mem[14'd7544] <= 32'hbdab4f91;
        mem[14'd7545] <= 32'hba8a0b7b;
        mem[14'd7546] <= 32'hbe10e579;
        mem[14'd7547] <= 32'h3dbc4861;
        mem[14'd7548] <= 32'h3e7aff02;
        mem[14'd7549] <= 32'h3ecc3e7c;
        mem[14'd7550] <= 32'h3cf962e2;
        mem[14'd7551] <= 32'h3e96fe4a;
        mem[14'd7552] <= 32'h3dfc1ba0;
        mem[14'd7553] <= 32'hbe2ca22c;
        mem[14'd7554] <= 32'hbcb3d515;
        mem[14'd7555] <= 32'h3d5f5b30;
        mem[14'd7556] <= 32'h3e1c25ff;
        mem[14'd7557] <= 32'hbc6d6471;
        mem[14'd7558] <= 32'h3daebea8;
        mem[14'd7559] <= 32'h3e04a599;
        mem[14'd7560] <= 32'h3da8a8e6;
        mem[14'd7561] <= 32'h3c365568;
        mem[14'd7562] <= 32'hbb88d372;
        mem[14'd7563] <= 32'hbb96d197;
        mem[14'd7564] <= 32'hbcdbac0a;
        mem[14'd7565] <= 32'hbc1ee830;
        mem[14'd7566] <= 32'h3c739fc5;
        mem[14'd7567] <= 32'hbc905a28;
        mem[14'd7568] <= 32'hbdbdbdbc;
        mem[14'd7569] <= 32'hbd9af74f;
        mem[14'd7570] <= 32'hbe183a1e;
        mem[14'd7571] <= 32'hbe9381e9;
        mem[14'd7572] <= 32'hbe93985c;
        mem[14'd7573] <= 32'hbe61106f;
        mem[14'd7574] <= 32'hbcee3236;
        mem[14'd7575] <= 32'h3e79aaba;
        mem[14'd7576] <= 32'h3e5e9185;
        mem[14'd7577] <= 32'h3eba681d;
        mem[14'd7578] <= 32'h3e6cd9f1;
        mem[14'd7579] <= 32'h3e1ec5c8;
        mem[14'd7580] <= 32'hbc16a36d;
        mem[14'd7581] <= 32'h3c81e8ed;
        mem[14'd7582] <= 32'hbd52f96d;
        mem[14'd7583] <= 32'hbd3adecc;
        mem[14'd7584] <= 32'hbe71d1a9;
        mem[14'd7585] <= 32'hbe556daf;
        mem[14'd7586] <= 32'hbe7bc02f;
        mem[14'd7587] <= 32'hbe4536be;
        mem[14'd7588] <= 32'hbde4964a;
        mem[14'd7589] <= 32'hbc2e24c1;
        mem[14'd7590] <= 32'hbb77645c;
        mem[14'd7591] <= 32'hbc5f8573;
        mem[14'd7592] <= 32'h395bd661;
        mem[14'd7593] <= 32'hbbc9b7e3;
        mem[14'd7594] <= 32'hbc351147;
        mem[14'd7595] <= 32'hbc1f9d37;
        mem[14'd7596] <= 32'hbdcf0ede;
        mem[14'd7597] <= 32'hbe5633e3;
        mem[14'd7598] <= 32'hbe7bd3ee;
        mem[14'd7599] <= 32'hbe761a67;
        mem[14'd7600] <= 32'hbe3bd605;
        mem[14'd7601] <= 32'hbd63c713;
        mem[14'd7602] <= 32'hbda3ffd0;
        mem[14'd7603] <= 32'hbd62a8e4;
        mem[14'd7604] <= 32'h3e4b89c0;
        mem[14'd7605] <= 32'h3ec3cd1d;
        mem[14'd7606] <= 32'h3ebb8968;
        mem[14'd7607] <= 32'h3db147cc;
        mem[14'd7608] <= 32'hbd74d6c9;
        mem[14'd7609] <= 32'hbdda9b1c;
        mem[14'd7610] <= 32'hbd83c8e3;
        mem[14'd7611] <= 32'hbe20d714;
        mem[14'd7612] <= 32'hbe9ff819;
        mem[14'd7613] <= 32'hbe9ce360;
        mem[14'd7614] <= 32'hbe6b7f8e;
        mem[14'd7615] <= 32'hbe7010d8;
        mem[14'd7616] <= 32'hbe317e12;
        mem[14'd7617] <= 32'hbcc94223;
        mem[14'd7618] <= 32'hbc87ca6c;
        mem[14'd7619] <= 32'hbad4cc56;
        mem[14'd7620] <= 32'h3c5c1687;
        mem[14'd7621] <= 32'h3c35959f;
        mem[14'd7622] <= 32'hbb5ac09d;
        mem[14'd7623] <= 32'h3b30b848;
        mem[14'd7624] <= 32'hbdf20d7b;
        mem[14'd7625] <= 32'hbe6c31dc;
        mem[14'd7626] <= 32'hbe29e406;
        mem[14'd7627] <= 32'hbd6927d0;
        mem[14'd7628] <= 32'h3d2d0171;
        mem[14'd7629] <= 32'h3d67027e;
        mem[14'd7630] <= 32'h3cdea419;
        mem[14'd7631] <= 32'h3d5bb864;
        mem[14'd7632] <= 32'h3ea3061c;
        mem[14'd7633] <= 32'h3e6cf62f;
        mem[14'd7634] <= 32'h3deabbf0;
        mem[14'd7635] <= 32'h3d810b92;
        mem[14'd7636] <= 32'h3df52e17;
        mem[14'd7637] <= 32'hbd0daee1;
        mem[14'd7638] <= 32'hbe6d10e7;
        mem[14'd7639] <= 32'hbeaebcf9;
        mem[14'd7640] <= 32'hbe9ed064;
        mem[14'd7641] <= 32'hbea98381;
        mem[14'd7642] <= 32'hbe941c0b;
        mem[14'd7643] <= 32'hbde6d166;
        mem[14'd7644] <= 32'hbe11bae8;
        mem[14'd7645] <= 32'hbd9dcedb;
        mem[14'd7646] <= 32'hbcd33f17;
        mem[14'd7647] <= 32'hbbc433b7;
        mem[14'd7648] <= 32'hbc155fb8;
        mem[14'd7649] <= 32'h3c59b63c;
        mem[14'd7650] <= 32'h3a679b01;
        mem[14'd7651] <= 32'hbd0d1dff;
        mem[14'd7652] <= 32'hbe044a4a;
        mem[14'd7653] <= 32'hbe4b82e4;
        mem[14'd7654] <= 32'hbdf5a82b;
        mem[14'd7655] <= 32'h3d9698b4;
        mem[14'd7656] <= 32'h3e130052;
        mem[14'd7657] <= 32'h3e68b2d4;
        mem[14'd7658] <= 32'h3dc6d520;
        mem[14'd7659] <= 32'h3e838087;
        mem[14'd7660] <= 32'h3ebc57bc;
        mem[14'd7661] <= 32'h3e41eade;
        mem[14'd7662] <= 32'h3d8f8532;
        mem[14'd7663] <= 32'hbdbd306d;
        mem[14'd7664] <= 32'h3dd3a611;
        mem[14'd7665] <= 32'hbdea6abe;
        mem[14'd7666] <= 32'hbe8a06ae;
        mem[14'd7667] <= 32'hbe2cc82e;
        mem[14'd7668] <= 32'hbdeb9f73;
        mem[14'd7669] <= 32'hbe109d4d;
        mem[14'd7670] <= 32'hbe0e1465;
        mem[14'd7671] <= 32'hbcb3bc94;
        mem[14'd7672] <= 32'hbd3d1022;
        mem[14'd7673] <= 32'hbe1180c1;
        mem[14'd7674] <= 32'hbcc41bb6;
        mem[14'd7675] <= 32'h3c36ab1f;
        mem[14'd7676] <= 32'h3c41cb67;
        mem[14'd7677] <= 32'hbc851431;
        mem[14'd7678] <= 32'h3b9797e5;
        mem[14'd7679] <= 32'hbd7f229f;
        mem[14'd7680] <= 32'hbe31b31c;
        mem[14'd7681] <= 32'hbdd3dcb4;
        mem[14'd7682] <= 32'h3c0c550c;
        mem[14'd7683] <= 32'h3d23b4c3;
        mem[14'd7684] <= 32'h3dde7831;
        mem[14'd7685] <= 32'h3e89632e;
        mem[14'd7686] <= 32'h3e85c57b;
        mem[14'd7687] <= 32'h3e82dbc7;
        mem[14'd7688] <= 32'h3e4bd87b;
        mem[14'd7689] <= 32'h3d7f3d68;
        mem[14'd7690] <= 32'hbe0294c5;
        mem[14'd7691] <= 32'hbd391500;
        mem[14'd7692] <= 32'hbdfd0a30;
        mem[14'd7693] <= 32'hbe3fa031;
        mem[14'd7694] <= 32'hbda38b35;
        mem[14'd7695] <= 32'hbd7668aa;
        mem[14'd7696] <= 32'hbb91faef;
        mem[14'd7697] <= 32'hbdee4f84;
        mem[14'd7698] <= 32'hbbccc705;
        mem[14'd7699] <= 32'h3d6cdbb8;
        mem[14'd7700] <= 32'hbd79b3ce;
        mem[14'd7701] <= 32'hbdf7dced;
        mem[14'd7702] <= 32'hbd01b61f;
        mem[14'd7703] <= 32'h3b1d3db2;
        mem[14'd7704] <= 32'hbc778548;
        mem[14'd7705] <= 32'hbb8c5cb9;
        mem[14'd7706] <= 32'h3b6637a1;
        mem[14'd7707] <= 32'hbdb93424;
        mem[14'd7708] <= 32'hbe4f7c8d;
        mem[14'd7709] <= 32'h3d65bf7f;
        mem[14'd7710] <= 32'h3db77f1b;
        mem[14'd7711] <= 32'hbab93fa5;
        mem[14'd7712] <= 32'h3d1918cd;
        mem[14'd7713] <= 32'h3e440804;
        mem[14'd7714] <= 32'h3e1ce615;
        mem[14'd7715] <= 32'hbda1a9a3;
        mem[14'd7716] <= 32'h3cd2e4cf;
        mem[14'd7717] <= 32'hbe03af79;
        mem[14'd7718] <= 32'hbe0c9ebc;
        mem[14'd7719] <= 32'hbd2f9da6;
        mem[14'd7720] <= 32'hbcdf95ee;
        mem[14'd7721] <= 32'hbbed03cf;
        mem[14'd7722] <= 32'h3d5e2c0e;
        mem[14'd7723] <= 32'h3cc80c0e;
        mem[14'd7724] <= 32'h3babee5d;
        mem[14'd7725] <= 32'hbb45ee0e;
        mem[14'd7726] <= 32'h3e357649;
        mem[14'd7727] <= 32'h3e065f5e;
        mem[14'd7728] <= 32'hbd646f17;
        mem[14'd7729] <= 32'hbdde3f43;
        mem[14'd7730] <= 32'h3adeaf36;
        mem[14'd7731] <= 32'hbc0f89ea;
        mem[14'd7732] <= 32'h3b7b842a;
        mem[14'd7733] <= 32'h3c9bffed;
        mem[14'd7734] <= 32'hbcb0ef6f;
        mem[14'd7735] <= 32'hbdf53bc5;
        mem[14'd7736] <= 32'hbe45cb39;
        mem[14'd7737] <= 32'h39a831a7;
        mem[14'd7738] <= 32'h3e0875a5;
        mem[14'd7739] <= 32'h3e860431;
        mem[14'd7740] <= 32'h3d91e67e;
        mem[14'd7741] <= 32'hbcdf6a84;
        mem[14'd7742] <= 32'h3ded12c6;
        mem[14'd7743] <= 32'hbe159881;
        mem[14'd7744] <= 32'h3d2d2b42;
        mem[14'd7745] <= 32'h3d0535c3;
        mem[14'd7746] <= 32'hbe0d3b7c;
        mem[14'd7747] <= 32'h3d5a080e;
        mem[14'd7748] <= 32'hbe2dbf9f;
        mem[14'd7749] <= 32'hbd821b7d;
        mem[14'd7750] <= 32'hbd09e926;
        mem[14'd7751] <= 32'hbc2d3998;
        mem[14'd7752] <= 32'h3dc104d1;
        mem[14'd7753] <= 32'h3e2d5e2a;
        mem[14'd7754] <= 32'h3e3a43fe;
        mem[14'd7755] <= 32'h3ddbe1cb;
        mem[14'd7756] <= 32'hbdb4e267;
        mem[14'd7757] <= 32'hbd83e0b0;
        mem[14'd7758] <= 32'hbc8eaa57;
        mem[14'd7759] <= 32'h3c204015;
        mem[14'd7760] <= 32'h3ba02d9d;
        mem[14'd7761] <= 32'hbb7c18bb;
        mem[14'd7762] <= 32'hbb6167b5;
        mem[14'd7763] <= 32'hbda1af00;
        mem[14'd7764] <= 32'hbdfc1041;
        mem[14'd7765] <= 32'hbd0a007b;
        mem[14'd7766] <= 32'h3e35e82b;
        mem[14'd7767] <= 32'h3e7d1131;
        mem[14'd7768] <= 32'h3ce9902b;
        mem[14'd7769] <= 32'h3dbcbece;
        mem[14'd7770] <= 32'hbd5ebaea;
        mem[14'd7771] <= 32'hbd710a23;
        mem[14'd7772] <= 32'hbdd03d3f;
        mem[14'd7773] <= 32'h3da47f10;
        mem[14'd7774] <= 32'hbc823cce;
        mem[14'd7775] <= 32'hbc9bf3e8;
        mem[14'd7776] <= 32'hbe038826;
        mem[14'd7777] <= 32'hbbe78979;
        mem[14'd7778] <= 32'hbd7d237b;
        mem[14'd7779] <= 32'hbd5d135d;
        mem[14'd7780] <= 32'h3dbde98d;
        mem[14'd7781] <= 32'h3d7f90ac;
        mem[14'd7782] <= 32'h3de7d403;
        mem[14'd7783] <= 32'h3b0352f2;
        mem[14'd7784] <= 32'hbdd9bf0b;
        mem[14'd7785] <= 32'hbcc3448f;
        mem[14'd7786] <= 32'hbc3b2e0b;
        mem[14'd7787] <= 32'hbc657dd7;
        mem[14'd7788] <= 32'hbaf71549;
        mem[14'd7789] <= 32'h3c6e9f7f;
        mem[14'd7790] <= 32'hbc27fecc;
        mem[14'd7791] <= 32'hbce7e164;
        mem[14'd7792] <= 32'hbdf7dad3;
        mem[14'd7793] <= 32'hbe1114c9;
        mem[14'd7794] <= 32'h3d4275ed;
        mem[14'd7795] <= 32'h3dfe0897;
        mem[14'd7796] <= 32'hbce17578;
        mem[14'd7797] <= 32'hbdbf17ed;
        mem[14'd7798] <= 32'hbbd7f5ad;
        mem[14'd7799] <= 32'h3de9173d;
        mem[14'd7800] <= 32'h3e11f855;
        mem[14'd7801] <= 32'h3e1e4f7c;
        mem[14'd7802] <= 32'h3e1bb3b8;
        mem[14'd7803] <= 32'h3d5a447a;
        mem[14'd7804] <= 32'hbd29cf3d;
        mem[14'd7805] <= 32'hbbea44c2;
        mem[14'd7806] <= 32'hbc4ea5ee;
        mem[14'd7807] <= 32'hbd84f944;
        mem[14'd7808] <= 32'hbca03c23;
        mem[14'd7809] <= 32'h3dafd04d;
        mem[14'd7810] <= 32'h3c9248db;
        mem[14'd7811] <= 32'hbccc243e;
        mem[14'd7812] <= 32'hbd1d1ce4;
        mem[14'd7813] <= 32'hbcb2b2db;
        mem[14'd7814] <= 32'hbbb883b4;
        mem[14'd7815] <= 32'h3bce83ad;
        mem[14'd7816] <= 32'hbc13ee64;
        mem[14'd7817] <= 32'hbc9855c4;
        mem[14'd7818] <= 32'h3c21513d;
        mem[14'd7819] <= 32'hbc3dcb8a;
        mem[14'd7820] <= 32'hbdd6b707;
        mem[14'd7821] <= 32'hbe98c3b0;
        mem[14'd7822] <= 32'hbe9e7c78;
        mem[14'd7823] <= 32'hbe30efa6;
        mem[14'd7824] <= 32'h3e002ff3;
        mem[14'd7825] <= 32'h3d6dd1fe;
        mem[14'd7826] <= 32'hbd0b5853;
        mem[14'd7827] <= 32'h3db1d27c;
        mem[14'd7828] <= 32'h3e487a08;
        mem[14'd7829] <= 32'h3eaf4fa7;
        mem[14'd7830] <= 32'h3e3bff45;
        mem[14'd7831] <= 32'h3e6ce046;
        mem[14'd7832] <= 32'h3e7dced3;
        mem[14'd7833] <= 32'h3dd17951;
        mem[14'd7834] <= 32'h3e0a1d40;
        mem[14'd7835] <= 32'h3e0aa45b;
        mem[14'd7836] <= 32'h3e01183a;
        mem[14'd7837] <= 32'h3da4a44d;
        mem[14'd7838] <= 32'hbc962538;
        mem[14'd7839] <= 32'h3ca01ef9;
        mem[14'd7840] <= 32'hbceb0d88;
        mem[14'd7841] <= 32'hbcb86f0c;
        mem[14'd7842] <= 32'hbc371933;
        mem[14'd7843] <= 32'h3a5e065d;
        mem[14'd7844] <= 32'hbc089dc3;
        mem[14'd7845] <= 32'h3c268586;
        mem[14'd7846] <= 32'hbbcd45ea;
        mem[14'd7847] <= 32'hbcc7c611;
        mem[14'd7848] <= 32'hbde53d41;
        mem[14'd7849] <= 32'hbe8ac0e6;
        mem[14'd7850] <= 32'hbea34f99;
        mem[14'd7851] <= 32'hbe8721a6;
        mem[14'd7852] <= 32'h3c9f0fe7;
        mem[14'd7853] <= 32'h3d853701;
        mem[14'd7854] <= 32'h3d9b0cd3;
        mem[14'd7855] <= 32'h3e548d6f;
        mem[14'd7856] <= 32'h3e5422d8;
        mem[14'd7857] <= 32'h3e0d13d5;
        mem[14'd7858] <= 32'h3e23ec29;
        mem[14'd7859] <= 32'h3e7a3219;
        mem[14'd7860] <= 32'h3eba1833;
        mem[14'd7861] <= 32'h3d1e4dca;
        mem[14'd7862] <= 32'h3e637765;
        mem[14'd7863] <= 32'h3ea38abe;
        mem[14'd7864] <= 32'h3dba4087;
        mem[14'd7865] <= 32'hbd5bc87f;
        mem[14'd7866] <= 32'hbd8a10fe;
        mem[14'd7867] <= 32'hbd3d0603;
        mem[14'd7868] <= 32'hbd1cef08;
        mem[14'd7869] <= 32'h3b440830;
        mem[14'd7870] <= 32'h3cba5643;
        mem[14'd7871] <= 32'hbc373515;
        mem[14'd7872] <= 32'hbae44fa7;
        mem[14'd7873] <= 32'hbbc58b5c;
        mem[14'd7874] <= 32'h3b8b5365;
        mem[14'd7875] <= 32'h3c51b792;
        mem[14'd7876] <= 32'hbd9b6a4c;
        mem[14'd7877] <= 32'hbe06152e;
        mem[14'd7878] <= 32'hbdf5c3ba;
        mem[14'd7879] <= 32'hbe1ffdc0;
        mem[14'd7880] <= 32'hbe484e7f;
        mem[14'd7881] <= 32'hbe41e499;
        mem[14'd7882] <= 32'hbd55a240;
        mem[14'd7883] <= 32'hbd08f6df;
        mem[14'd7884] <= 32'hbd986fb7;
        mem[14'd7885] <= 32'hbd77668a;
        mem[14'd7886] <= 32'h3db90e58;
        mem[14'd7887] <= 32'h3e1e1a37;
        mem[14'd7888] <= 32'h3e13e89d;
        mem[14'd7889] <= 32'h3e11eeec;
        mem[14'd7890] <= 32'h3dad147b;
        mem[14'd7891] <= 32'h3d72f011;
        mem[14'd7892] <= 32'h3be405ab;
        mem[14'd7893] <= 32'hbd042d3f;
        mem[14'd7894] <= 32'hbcfce3f1;
        mem[14'd7895] <= 32'hbcbd1ebc;
        mem[14'd7896] <= 32'hbb756e8e;
        mem[14'd7897] <= 32'hbb9b670c;
        mem[14'd7898] <= 32'h3b6f7cd5;
        mem[14'd7899] <= 32'hbba930fd;
        mem[14'd7900] <= 32'h3b7cd567;
        mem[14'd7901] <= 32'hbc182767;
        mem[14'd7902] <= 32'h3c0b32d9;
        mem[14'd7903] <= 32'hbb60c0d2;
        mem[14'd7904] <= 32'hbc9447bd;
        mem[14'd7905] <= 32'hbc864bf4;
        mem[14'd7906] <= 32'hbca0ed34;
        mem[14'd7907] <= 32'hbc436029;
        mem[14'd7908] <= 32'hbcac342c;
        mem[14'd7909] <= 32'hbd63c830;
        mem[14'd7910] <= 32'hbd9f23c3;
        mem[14'd7911] <= 32'hbdadaeb9;
        mem[14'd7912] <= 32'hbdaf8845;
        mem[14'd7913] <= 32'hbdb48f00;
        mem[14'd7914] <= 32'hbdc7e7ac;
        mem[14'd7915] <= 32'hbdd2b784;
        mem[14'd7916] <= 32'hbdb91aa2;
        mem[14'd7917] <= 32'hbd517f5d;
        mem[14'd7918] <= 32'hbcc35ba6;
        mem[14'd7919] <= 32'hbcf77905;
        mem[14'd7920] <= 32'hbcfb7844;
        mem[14'd7921] <= 32'hbc890094;
        mem[14'd7922] <= 32'hbc67ca3f;
        mem[14'd7923] <= 32'hbc7caac7;
        mem[14'd7924] <= 32'hba5e22df;
        mem[14'd7925] <= 32'hbc627191;
        mem[14'd7926] <= 32'h3c922d9e;
        mem[14'd7927] <= 32'hbc2f46dc;
        mem[14'd7928] <= 32'hbb520dec;
        mem[14'd7929] <= 32'hbb38f301;
        mem[14'd7930] <= 32'h3bc7ac6d;
        mem[14'd7931] <= 32'hbc443ca2;
        mem[14'd7932] <= 32'h3c2632b8;
        mem[14'd7933] <= 32'hbc10f9c4;
        mem[14'd7934] <= 32'h3a02eaaf;
        mem[14'd7935] <= 32'h3bbc8fef;
        mem[14'd7936] <= 32'h3c50ba66;
        mem[14'd7937] <= 32'hbc538458;
        mem[14'd7938] <= 32'h3c12ddab;
        mem[14'd7939] <= 32'h3bd020e3;
        mem[14'd7940] <= 32'hbbfd9850;
        mem[14'd7941] <= 32'hbad68225;
        mem[14'd7942] <= 32'hbb8f3cdb;
        mem[14'd7943] <= 32'hba78e7c9;
        mem[14'd7944] <= 32'hbbce2836;
        mem[14'd7945] <= 32'hba8e7408;
        mem[14'd7946] <= 32'hbc9acb64;
        mem[14'd7947] <= 32'h3c35ac6a;
        mem[14'd7948] <= 32'hbc3f0466;
        mem[14'd7949] <= 32'hbc86f62e;
        mem[14'd7950] <= 32'hbaeb7b20;
        mem[14'd7951] <= 32'h3c2f2a36;
        mem[14'd7952] <= 32'hbb92b032;
        mem[14'd7953] <= 32'h3c4cf646;
        mem[14'd7954] <= 32'hbbdf7527;
        mem[14'd7955] <= 32'h3bdf4ba5;
        mem[14'd7956] <= 32'hbbd0d48a;
        mem[14'd7957] <= 32'h3b14ac73;
        mem[14'd7958] <= 32'hbc2df121;
        mem[14'd7959] <= 32'h3c95fd69;
        mem[14'd7960] <= 32'hbb32b5c0;
        mem[14'd7961] <= 32'h3c002d11;
        mem[14'd7962] <= 32'h3c3d74d7;
        mem[14'd7963] <= 32'hba066963;
        mem[14'd7964] <= 32'h3c1cb750;
        mem[14'd7965] <= 32'h3bba7e84;
        mem[14'd7966] <= 32'hbc12077b;
        mem[14'd7967] <= 32'hbc2a3b0f;
        mem[14'd7968] <= 32'hbb2d4bec;
        mem[14'd7969] <= 32'h3c4c9c03;
        mem[14'd7970] <= 32'h3c01a473;
        mem[14'd7971] <= 32'hbae9dbc0;
        mem[14'd7972] <= 32'hbc7b96fd;
        mem[14'd7973] <= 32'h3a96c846;
        mem[14'd7974] <= 32'h3c04452a;
        mem[14'd7975] <= 32'hbc307a59;
        mem[14'd7976] <= 32'hbc7b6f18;
        mem[14'd7977] <= 32'h3c309a4d;
        mem[14'd7978] <= 32'hbac0eeed;
        mem[14'd7979] <= 32'hbc86c607;
        mem[14'd7980] <= 32'h3bae77c7;
        mem[14'd7981] <= 32'hbbe41492;
        mem[14'd7982] <= 32'h3c0af875;
        mem[14'd7983] <= 32'h3c2ccc45;
        mem[14'd7984] <= 32'h3a73e543;
        mem[14'd7985] <= 32'hbbc81740;
        mem[14'd7986] <= 32'hbbff0a9c;
        mem[14'd7987] <= 32'hbb747c61;
        mem[14'd7988] <= 32'h3cc1ebd7;
        mem[14'd7989] <= 32'hbc825dbd;
        mem[14'd7990] <= 32'h3c5f7f03;
        mem[14'd7991] <= 32'hbcc4f047;
        mem[14'd7992] <= 32'h3c8b6744;
        mem[14'd7993] <= 32'h3c821ea6;
        mem[14'd7994] <= 32'h3bf2e05b;
        mem[14'd7995] <= 32'hbb6f6442;
        mem[14'd7996] <= 32'h3be642c6;
        mem[14'd7997] <= 32'h3985e9f9;
        mem[14'd7998] <= 32'hbaf4f499;
        mem[14'd7999] <= 32'hbc168c74;
        mem[14'd8000] <= 32'hbc4e70ac;
        mem[14'd8001] <= 32'hbb8bf0ad;
        mem[14'd8002] <= 32'hbbcff39b;
        mem[14'd8003] <= 32'h3bf48a97;
        mem[14'd8004] <= 32'h3b180435;
        mem[14'd8005] <= 32'h3c0d40f2;
        mem[14'd8006] <= 32'hbb6ac026;
        mem[14'd8007] <= 32'h39fe145e;
        mem[14'd8008] <= 32'h3c5c75dd;
        mem[14'd8009] <= 32'hb72ccb96;
        mem[14'd8010] <= 32'h3c801b34;
        mem[14'd8011] <= 32'h3cb7b6bb;
        mem[14'd8012] <= 32'h3ad9b2e4;
        mem[14'd8013] <= 32'hbaaee3e5;
        mem[14'd8014] <= 32'hbc0117a3;
        mem[14'd8015] <= 32'h3ccd10c6;
        mem[14'd8016] <= 32'hbb28e4d7;
        mem[14'd8017] <= 32'h3ca903b6;
        mem[14'd8018] <= 32'h3b8880d5;
        mem[14'd8019] <= 32'h3be22254;
        mem[14'd8020] <= 32'hbb1abe17;
        mem[14'd8021] <= 32'hbbdd7811;
        mem[14'd8022] <= 32'hbad6dfa1;
        mem[14'd8023] <= 32'h3b0ddb19;
        mem[14'd8024] <= 32'hbcc6be04;
        mem[14'd8025] <= 32'hbcc1b830;
        mem[14'd8026] <= 32'hbd0b329d;
        mem[14'd8027] <= 32'hbd1b2199;
        mem[14'd8028] <= 32'hbd038b41;
        mem[14'd8029] <= 32'hbc9d6e33;
        mem[14'd8030] <= 32'hbcc85e86;
        mem[14'd8031] <= 32'hbc8529c9;
        mem[14'd8032] <= 32'h3ac95a44;
        mem[14'd8033] <= 32'h3c1efb4a;
        mem[14'd8034] <= 32'hba467390;
        mem[14'd8035] <= 32'hbc005b1a;
        mem[14'd8036] <= 32'h3bba13a8;
        mem[14'd8037] <= 32'hbc426ddf;
        mem[14'd8038] <= 32'hbb3563be;
        mem[14'd8039] <= 32'hbb709ad9;
        mem[14'd8040] <= 32'h3ca1d02a;
        mem[14'd8041] <= 32'hbb0c1c46;
        mem[14'd8042] <= 32'h3cf30211;
        mem[14'd8043] <= 32'hbb8f3a43;
        mem[14'd8044] <= 32'hbb608a8f;
        mem[14'd8045] <= 32'h3c13656d;
        mem[14'd8046] <= 32'h390db3ab;
        mem[14'd8047] <= 32'h3b812d79;
        mem[14'd8048] <= 32'hbbc6b3c4;
        mem[14'd8049] <= 32'hbb32dfc2;
        mem[14'd8050] <= 32'hbcdbf364;
        mem[14'd8051] <= 32'hbd5c6bba;
        mem[14'd8052] <= 32'hbd93e4e1;
        mem[14'd8053] <= 32'hbdbd44f0;
        mem[14'd8054] <= 32'hbdd5bc48;
        mem[14'd8055] <= 32'hbe1ca673;
        mem[14'd8056] <= 32'hbdc9328d;
        mem[14'd8057] <= 32'hbdc11a32;
        mem[14'd8058] <= 32'hbd29db95;
        mem[14'd8059] <= 32'hbd235a4e;
        mem[14'd8060] <= 32'hbd6c7510;
        mem[14'd8061] <= 32'hbc6282e2;
        mem[14'd8062] <= 32'hbb810743;
        mem[14'd8063] <= 32'hbc2cf4fc;
        mem[14'd8064] <= 32'h3c80d549;
        mem[14'd8065] <= 32'h3c0f73c0;
        mem[14'd8066] <= 32'hbbac9c6f;
        mem[14'd8067] <= 32'hbae41102;
        mem[14'd8068] <= 32'hbaaf6a29;
        mem[14'd8069] <= 32'h3b1fed51;
        mem[14'd8070] <= 32'h3c267cc8;
        mem[14'd8071] <= 32'hb9e6590b;
        mem[14'd8072] <= 32'h3bd28576;
        mem[14'd8073] <= 32'h3c26bde8;
        mem[14'd8074] <= 32'hbc4b9d6b;
        mem[14'd8075] <= 32'hbcc19a73;
        mem[14'd8076] <= 32'hbd746afc;
        mem[14'd8077] <= 32'hbd95620a;
        mem[14'd8078] <= 32'hbdd4e390;
        mem[14'd8079] <= 32'hbe111a08;
        mem[14'd8080] <= 32'hbe43fe2a;
        mem[14'd8081] <= 32'hbe67e4bf;
        mem[14'd8082] <= 32'hbe9015a6;
        mem[14'd8083] <= 32'hbea22f9a;
        mem[14'd8084] <= 32'hbeab91c6;
        mem[14'd8085] <= 32'hbe9034a9;
        mem[14'd8086] <= 32'hbe54eeed;
        mem[14'd8087] <= 32'hbe49bb5d;
        mem[14'd8088] <= 32'hbe1248a1;
        mem[14'd8089] <= 32'hbdda391d;
        mem[14'd8090] <= 32'hbd894531;
        mem[14'd8091] <= 32'hbd140565;
        mem[14'd8092] <= 32'h3a985743;
        mem[14'd8093] <= 32'h3be97095;
        mem[14'd8094] <= 32'hba5f22bc;
        mem[14'd8095] <= 32'h3c5ba4a0;
        mem[14'd8096] <= 32'hbcacf5ea;
        mem[14'd8097] <= 32'hbad9d88f;
        mem[14'd8098] <= 32'hbb89c018;
        mem[14'd8099] <= 32'h3c6b7e32;
        mem[14'd8100] <= 32'h3bfa25d7;
        mem[14'd8101] <= 32'hbc663c9e;
        mem[14'd8102] <= 32'hbd3e4f36;
        mem[14'd8103] <= 32'hbdbfd911;
        mem[14'd8104] <= 32'hbe0d8ef5;
        mem[14'd8105] <= 32'hbe3a0a8b;
        mem[14'd8106] <= 32'hbdf40af0;
        mem[14'd8107] <= 32'h3db65842;
        mem[14'd8108] <= 32'h3db6b74b;
        mem[14'd8109] <= 32'h3de3ac07;
        mem[14'd8110] <= 32'hbda0e367;
        mem[14'd8111] <= 32'hbdc030e3;
        mem[14'd8112] <= 32'hbea542c8;
        mem[14'd8113] <= 32'hbe8ec778;
        mem[14'd8114] <= 32'hbe8f1507;
        mem[14'd8115] <= 32'hbe6a9144;
        mem[14'd8116] <= 32'hbe7c6b3e;
        mem[14'd8117] <= 32'hbe744f3d;
        mem[14'd8118] <= 32'hbe63e5c5;
        mem[14'd8119] <= 32'hbe07a312;
        mem[14'd8120] <= 32'hbd92a705;
        mem[14'd8121] <= 32'hbcaa7e2c;
        mem[14'd8122] <= 32'hbc6fe4e4;
        mem[14'd8123] <= 32'h3c9ed68c;
        mem[14'd8124] <= 32'hbc73b4e2;
        mem[14'd8125] <= 32'hbbb3498c;
        mem[14'd8126] <= 32'hbc5fa592;
        mem[14'd8127] <= 32'hbca2f809;
        mem[14'd8128] <= 32'hbd28e964;
        mem[14'd8129] <= 32'hbe1b72e3;
        mem[14'd8130] <= 32'hbe4c19b0;
        mem[14'd8131] <= 32'hbe6eaa94;
        mem[14'd8132] <= 32'hbe5829fa;
        mem[14'd8133] <= 32'hbdcc3627;
        mem[14'd8134] <= 32'hbca8e47f;
        mem[14'd8135] <= 32'h3e060f58;
        mem[14'd8136] <= 32'h3dfcf089;
        mem[14'd8137] <= 32'h3e8c2cf6;
        mem[14'd8138] <= 32'h3e8e28f9;
        mem[14'd8139] <= 32'h3e565f45;
        mem[14'd8140] <= 32'h3e780488;
        mem[14'd8141] <= 32'h3e654eca;
        mem[14'd8142] <= 32'h3e4dd782;
        mem[14'd8143] <= 32'h3c341f86;
        mem[14'd8144] <= 32'hbc5218a7;
        mem[14'd8145] <= 32'hbe1e7f09;
        mem[14'd8146] <= 32'hbe89c3da;
        mem[14'd8147] <= 32'hbe8373df;
        mem[14'd8148] <= 32'hbe13c4f2;
        mem[14'd8149] <= 32'hbd8e591b;
        mem[14'd8150] <= 32'hbc968e53;
        mem[14'd8151] <= 32'hbcaec9e2;
        mem[14'd8152] <= 32'hbc380fbf;
        mem[14'd8153] <= 32'hbbebad95;
        mem[14'd8154] <= 32'hbc9b25f1;
        mem[14'd8155] <= 32'hbd39ecc3;
        mem[14'd8156] <= 32'hbe015b8d;
        mem[14'd8157] <= 32'hbe8855cc;
        mem[14'd8158] <= 32'hbe7adadb;
        mem[14'd8159] <= 32'hbe9555e0;
        mem[14'd8160] <= 32'hbdc74a2a;
        mem[14'd8161] <= 32'h3bb9e76b;
        mem[14'd8162] <= 32'h3d58e4fa;
        mem[14'd8163] <= 32'h3da5d6ee;
        mem[14'd8164] <= 32'h3e943649;
        mem[14'd8165] <= 32'h3ed82fdf;
        mem[14'd8166] <= 32'h3efe30ed;
        mem[14'd8167] <= 32'h3f071a09;
        mem[14'd8168] <= 32'h3efef13d;
        mem[14'd8169] <= 32'h3e9326fe;
        mem[14'd8170] <= 32'h3e2a3d36;
        mem[14'd8171] <= 32'h3daaed30;
        mem[14'd8172] <= 32'h3db4cd5a;
        mem[14'd8173] <= 32'hbb885b51;
        mem[14'd8174] <= 32'hbe3fb281;
        mem[14'd8175] <= 32'hbe7a765a;
        mem[14'd8176] <= 32'hbe56b56d;
        mem[14'd8177] <= 32'hbdba8c0d;
        mem[14'd8178] <= 32'hbd16ecb4;
        mem[14'd8179] <= 32'hbb850fa9;
        mem[14'd8180] <= 32'hbc793f46;
        mem[14'd8181] <= 32'hbcf522ef;
        mem[14'd8182] <= 32'hbd074779;
        mem[14'd8183] <= 32'hbdf4efe3;
        mem[14'd8184] <= 32'hbe4da994;
        mem[14'd8185] <= 32'hbe775c3d;
        mem[14'd8186] <= 32'hbe04d5c2;
        mem[14'd8187] <= 32'hbe38f3fc;
        mem[14'd8188] <= 32'h3da972de;
        mem[14'd8189] <= 32'hbd42f508;
        mem[14'd8190] <= 32'hbce6060d;
        mem[14'd8191] <= 32'hbd8bd2e1;
        mem[14'd8192] <= 32'hbe25833d;
        mem[14'd8193] <= 32'h3e099a48;
        mem[14'd8194] <= 32'h3ea18752;
        mem[14'd8195] <= 32'h3e5dbd8d;
        mem[14'd8196] <= 32'h3e275faf;
        mem[14'd8197] <= 32'h3d17f7b0;
        mem[14'd8198] <= 32'h3d7ba405;
        mem[14'd8199] <= 32'hbb654e2f;
        mem[14'd8200] <= 32'hbd26d0c7;
        mem[14'd8201] <= 32'h3dfa3fac;
        mem[14'd8202] <= 32'hbdbfedaf;
        mem[14'd8203] <= 32'hbe489130;
        mem[14'd8204] <= 32'hbe4245a3;
        mem[14'd8205] <= 32'hbde50c8f;
        mem[14'd8206] <= 32'hbcc9bc63;
        mem[14'd8207] <= 32'hbbc330d2;
        mem[14'd8208] <= 32'h3c1db4f6;
        mem[14'd8209] <= 32'hbcd5022d;
        mem[14'd8210] <= 32'hbd88dd7b;
        mem[14'd8211] <= 32'hbe1d9f51;
        mem[14'd8212] <= 32'hbe6c9fbe;
        mem[14'd8213] <= 32'hbde3c483;
        mem[14'd8214] <= 32'h3dbf90b9;
        mem[14'd8215] <= 32'h39611b6e;
        mem[14'd8216] <= 32'h3d361856;
        mem[14'd8217] <= 32'h3beb2448;
        mem[14'd8218] <= 32'h3dfc4987;
        mem[14'd8219] <= 32'h3d2e2c68;
        mem[14'd8220] <= 32'h3b18b20e;
        mem[14'd8221] <= 32'h3d7ea975;
        mem[14'd8222] <= 32'h3e4ac675;
        mem[14'd8223] <= 32'h3e81ff42;
        mem[14'd8224] <= 32'hbb1b3ee7;
        mem[14'd8225] <= 32'hba6ae6cf;
        mem[14'd8226] <= 32'h3db0a531;
        mem[14'd8227] <= 32'h3beec8dc;
        mem[14'd8228] <= 32'h3c983ce1;
        mem[14'd8229] <= 32'hbe01ae0f;
        mem[14'd8230] <= 32'hbe0236f8;
        mem[14'd8231] <= 32'hbe532cd6;
        mem[14'd8232] <= 32'hbe395278;
        mem[14'd8233] <= 32'hbddbe5a2;
        mem[14'd8234] <= 32'hbcd03b2c;
        mem[14'd8235] <= 32'h3c65266c;
        mem[14'd8236] <= 32'hba519b95;
        mem[14'd8237] <= 32'hbcbeb6cf;
        mem[14'd8238] <= 32'hbd76d02a;
        mem[14'd8239] <= 32'hbe12b167;
        mem[14'd8240] <= 32'hbe37d492;
        mem[14'd8241] <= 32'h3d02128b;
        mem[14'd8242] <= 32'h3e4abbf2;
        mem[14'd8243] <= 32'h3d6cd557;
        mem[14'd8244] <= 32'h3e2677bf;
        mem[14'd8245] <= 32'h3dbb7876;
        mem[14'd8246] <= 32'h3e126207;
        mem[14'd8247] <= 32'h3e4ee1fc;
        mem[14'd8248] <= 32'h3e07ab18;
        mem[14'd8249] <= 32'hbe1c345e;
        mem[14'd8250] <= 32'hbc17c832;
        mem[14'd8251] <= 32'hbd4ff811;
        mem[14'd8252] <= 32'h3c340185;
        mem[14'd8253] <= 32'h3b4298c7;
        mem[14'd8254] <= 32'h3d80686c;
        mem[14'd8255] <= 32'h3c7552a7;
        mem[14'd8256] <= 32'h3ce780a7;
        mem[14'd8257] <= 32'hbac2ddf5;
        mem[14'd8258] <= 32'hbd037b2c;
        mem[14'd8259] <= 32'hbdfd9b4e;
        mem[14'd8260] <= 32'hbe4ac2c5;
        mem[14'd8261] <= 32'hbdbc994c;
        mem[14'd8262] <= 32'hbd0f4a06;
        mem[14'd8263] <= 32'hbba1403a;
        mem[14'd8264] <= 32'hbb1fe953;
        mem[14'd8265] <= 32'hbd28620f;
        mem[14'd8266] <= 32'hbdf39e78;
        mem[14'd8267] <= 32'hbe276f04;
        mem[14'd8268] <= 32'hbcd810cf;
        mem[14'd8269] <= 32'h3e6caa8a;
        mem[14'd8270] <= 32'h3e80a750;
        mem[14'd8271] <= 32'h3e26889c;
        mem[14'd8272] <= 32'h3ec5bf70;
        mem[14'd8273] <= 32'h3e52bc69;
        mem[14'd8274] <= 32'h3e80d089;
        mem[14'd8275] <= 32'h3e99c9d2;
        mem[14'd8276] <= 32'h3d7bdf5b;
        mem[14'd8277] <= 32'hbce06d47;
        mem[14'd8278] <= 32'h3d137ca9;
        mem[14'd8279] <= 32'h3e392c09;
        mem[14'd8280] <= 32'h3e7e1c4f;
        mem[14'd8281] <= 32'h3eafdb8c;
        mem[14'd8282] <= 32'h3e6af7e3;
        mem[14'd8283] <= 32'h3e3ed7fe;
        mem[14'd8284] <= 32'h3edf1f8e;
        mem[14'd8285] <= 32'h3e9b989f;
        mem[14'd8286] <= 32'h3e5a7774;
        mem[14'd8287] <= 32'hbc8c7bd4;
        mem[14'd8288] <= 32'hbe1c0b15;
        mem[14'd8289] <= 32'hbd84f36e;
        mem[14'd8290] <= 32'hbbc757d0;
        mem[14'd8291] <= 32'h3c8727f0;
        mem[14'd8292] <= 32'h3a96b28d;
        mem[14'd8293] <= 32'hbcac7e85;
        mem[14'd8294] <= 32'hbda3c432;
        mem[14'd8295] <= 32'hbdebe79a;
        mem[14'd8296] <= 32'h3e2a384e;
        mem[14'd8297] <= 32'h3eb2acbf;
        mem[14'd8298] <= 32'h3ea284eb;
        mem[14'd8299] <= 32'h3e3986c5;
        mem[14'd8300] <= 32'h3e629420;
        mem[14'd8301] <= 32'h3e8fb2c8;
        mem[14'd8302] <= 32'h3e7eb7ad;
        mem[14'd8303] <= 32'h3e14a1ee;
        mem[14'd8304] <= 32'hbe53b84f;
        mem[14'd8305] <= 32'h3cd2c66b;
        mem[14'd8306] <= 32'h3e7a8476;
        mem[14'd8307] <= 32'h3e9528d4;
        mem[14'd8308] <= 32'h3e95a909;
        mem[14'd8309] <= 32'h3eb45cd0;
        mem[14'd8310] <= 32'h3ea75d9f;
        mem[14'd8311] <= 32'h3eca6391;
        mem[14'd8312] <= 32'h3eb9fb16;
        mem[14'd8313] <= 32'h3ec8184f;
        mem[14'd8314] <= 32'h3e84f297;
        mem[14'd8315] <= 32'h3dd93d58;
        mem[14'd8316] <= 32'hbe0b13a1;
        mem[14'd8317] <= 32'hbda0644c;
        mem[14'd8318] <= 32'hbc78c00b;
        mem[14'd8319] <= 32'h3c8ab134;
        mem[14'd8320] <= 32'hbc80f360;
        mem[14'd8321] <= 32'hbb3b7dfa;
        mem[14'd8322] <= 32'hbd8f3a33;
        mem[14'd8323] <= 32'hbd2e2a3a;
        mem[14'd8324] <= 32'h3ea7456f;
        mem[14'd8325] <= 32'h3eacab2d;
        mem[14'd8326] <= 32'h3e2f9147;
        mem[14'd8327] <= 32'h3e5ec43a;
        mem[14'd8328] <= 32'h3e5332ac;
        mem[14'd8329] <= 32'h3d908029;
        mem[14'd8330] <= 32'h3de92248;
        mem[14'd8331] <= 32'hbd1203ed;
        mem[14'd8332] <= 32'hbe4f06ec;
        mem[14'd8333] <= 32'h3dbcb810;
        mem[14'd8334] <= 32'h3e690637;
        mem[14'd8335] <= 32'h3e870e68;
        mem[14'd8336] <= 32'h3ec3af05;
        mem[14'd8337] <= 32'h3e9dbb18;
        mem[14'd8338] <= 32'h3e80da9a;
        mem[14'd8339] <= 32'h3ecc3af5;
        mem[14'd8340] <= 32'h3ea22f81;
        mem[14'd8341] <= 32'h3eac6a31;
        mem[14'd8342] <= 32'h3dcaae60;
        mem[14'd8343] <= 32'hbe25a42a;
        mem[14'd8344] <= 32'hbe630ef8;
        mem[14'd8345] <= 32'hbddef03f;
        mem[14'd8346] <= 32'hbceb985b;
        mem[14'd8347] <= 32'hbbb3e6ca;
        mem[14'd8348] <= 32'hbc9dd570;
        mem[14'd8349] <= 32'h3bf455fc;
        mem[14'd8350] <= 32'hbd0a0979;
        mem[14'd8351] <= 32'h3cb8f201;
        mem[14'd8352] <= 32'h3e5aefb9;
        mem[14'd8353] <= 32'h3e07b271;
        mem[14'd8354] <= 32'h3e316015;
        mem[14'd8355] <= 32'h3e0a52f3;
        mem[14'd8356] <= 32'h3d5e9729;
        mem[14'd8357] <= 32'h3bad98f9;
        mem[14'd8358] <= 32'h3d05c3cb;
        mem[14'd8359] <= 32'hbd254b26;
        mem[14'd8360] <= 32'hbdb402d2;
        mem[14'd8361] <= 32'h3d818205;
        mem[14'd8362] <= 32'h3cd80dd4;
        mem[14'd8363] <= 32'h3e4bf102;
        mem[14'd8364] <= 32'h3eab38bc;
        mem[14'd8365] <= 32'h3e92077f;
        mem[14'd8366] <= 32'h3e32589f;
        mem[14'd8367] <= 32'h3dd263c8;
        mem[14'd8368] <= 32'h3e4206af;
        mem[14'd8369] <= 32'h3e0a8898;
        mem[14'd8370] <= 32'hbd8b778d;
        mem[14'd8371] <= 32'hbe9dc558;
        mem[14'd8372] <= 32'hbe89489c;
        mem[14'd8373] <= 32'hbdb988a9;
        mem[14'd8374] <= 32'hbc90ccc2;
        mem[14'd8375] <= 32'h3c457cde;
        mem[14'd8376] <= 32'h3b78f49a;
        mem[14'd8377] <= 32'h3bd38618;
        mem[14'd8378] <= 32'hbd05e103;
        mem[14'd8379] <= 32'hbcd4b278;
        mem[14'd8380] <= 32'h3db430b7;
        mem[14'd8381] <= 32'h3da5ebfa;
        mem[14'd8382] <= 32'h3d33b51d;
        mem[14'd8383] <= 32'h3d2bf372;
        mem[14'd8384] <= 32'h3d850a84;
        mem[14'd8385] <= 32'hbdbcf0e4;
        mem[14'd8386] <= 32'h3d484ff0;
        mem[14'd8387] <= 32'h3d235c9e;
        mem[14'd8388] <= 32'hbd7fbbdb;
        mem[14'd8389] <= 32'hbdee8a91;
        mem[14'd8390] <= 32'hbe368ee5;
        mem[14'd8391] <= 32'h3e10e948;
        mem[14'd8392] <= 32'h3ea2d619;
        mem[14'd8393] <= 32'h3ea34c2a;
        mem[14'd8394] <= 32'h3df6e2b0;
        mem[14'd8395] <= 32'h3d21496f;
        mem[14'd8396] <= 32'h3d2aa717;
        mem[14'd8397] <= 32'hbdbb6cff;
        mem[14'd8398] <= 32'hbe634490;
        mem[14'd8399] <= 32'hbea659cb;
        mem[14'd8400] <= 32'hbe74ecd8;
        mem[14'd8401] <= 32'hbd4cb11b;
        mem[14'd8402] <= 32'hbc4e0bde;
        mem[14'd8403] <= 32'hbc6624ca;
        mem[14'd8404] <= 32'hbbfdc676;
        mem[14'd8405] <= 32'hbbd4fbe6;
        mem[14'd8406] <= 32'hbd1b9622;
        mem[14'd8407] <= 32'hbd1dd67f;
        mem[14'd8408] <= 32'h3d20b82e;
        mem[14'd8409] <= 32'h3c9ab1ea;
        mem[14'd8410] <= 32'hbdb01c79;
        mem[14'd8411] <= 32'hbcab175e;
        mem[14'd8412] <= 32'h3de236b6;
        mem[14'd8413] <= 32'hbdc4082e;
        mem[14'd8414] <= 32'h3d0863e5;
        mem[14'd8415] <= 32'h3d85f87a;
        mem[14'd8416] <= 32'hbd97e8dc;
        mem[14'd8417] <= 32'hbe635f23;
        mem[14'd8418] <= 32'hbde960ee;
        mem[14'd8419] <= 32'h3d01e532;
        mem[14'd8420] <= 32'h3e6ed78d;
        mem[14'd8421] <= 32'h3e4cf552;
        mem[14'd8422] <= 32'h3d47e038;
        mem[14'd8423] <= 32'hbe1886fc;
        mem[14'd8424] <= 32'hbe1a878e;
        mem[14'd8425] <= 32'hbe858a15;
        mem[14'd8426] <= 32'hbe64bd02;
        mem[14'd8427] <= 32'hbeb7054c;
        mem[14'd8428] <= 32'hbe8709f3;
        mem[14'd8429] <= 32'hbd9df454;
        mem[14'd8430] <= 32'hbd07c9b7;
        mem[14'd8431] <= 32'hbbc4c1f2;
        mem[14'd8432] <= 32'h3ae68502;
        mem[14'd8433] <= 32'hbad969f7;
        mem[14'd8434] <= 32'hbca3bbb7;
        mem[14'd8435] <= 32'hbd761fb1;
        mem[14'd8436] <= 32'hbe10da1b;
        mem[14'd8437] <= 32'hbe25bc62;
        mem[14'd8438] <= 32'hbe16eb31;
        mem[14'd8439] <= 32'h3b9c2af5;
        mem[14'd8440] <= 32'h3d70a31e;
        mem[14'd8441] <= 32'hbcb91a4b;
        mem[14'd8442] <= 32'h3d8282b8;
        mem[14'd8443] <= 32'h3c88faf8;
        mem[14'd8444] <= 32'h3c318f64;
        mem[14'd8445] <= 32'hbd09cefc;
        mem[14'd8446] <= 32'hbd6e1856;
        mem[14'd8447] <= 32'h3e689e55;
        mem[14'd8448] <= 32'h3d1d1d57;
        mem[14'd8449] <= 32'h3d4f4400;
        mem[14'd8450] <= 32'hbd3c2fb8;
        mem[14'd8451] <= 32'hbdf887ec;
        mem[14'd8452] <= 32'hbe08c1f7;
        mem[14'd8453] <= 32'hbe730779;
        mem[14'd8454] <= 32'hbe9dfb7b;
        mem[14'd8455] <= 32'hbeb025d7;
        mem[14'd8456] <= 32'hbe85de92;
        mem[14'd8457] <= 32'hbd51710c;
        mem[14'd8458] <= 32'hbc0a0142;
        mem[14'd8459] <= 32'hbb4ffd9b;
        mem[14'd8460] <= 32'hbc162b09;
        mem[14'd8461] <= 32'hbbaa7e60;
        mem[14'd8462] <= 32'hb9cb71b7;
        mem[14'd8463] <= 32'hbdee45ba;
        mem[14'd8464] <= 32'hbe3025b6;
        mem[14'd8465] <= 32'hbe7e83bf;
        mem[14'd8466] <= 32'hbdfe7048;
        mem[14'd8467] <= 32'hbdbf4984;
        mem[14'd8468] <= 32'hbdde8fbd;
        mem[14'd8469] <= 32'hbcc2d09f;
        mem[14'd8470] <= 32'h3e1bef2a;
        mem[14'd8471] <= 32'h3da2b833;
        mem[14'd8472] <= 32'hbe4e4e76;
        mem[14'd8473] <= 32'hbe29430a;
        mem[14'd8474] <= 32'h3dd44e73;
        mem[14'd8475] <= 32'h3de25001;
        mem[14'd8476] <= 32'hbdd2a3c7;
        mem[14'd8477] <= 32'hbda1d35c;
        mem[14'd8478] <= 32'hbe19c7ae;
        mem[14'd8479] <= 32'hbd6f2a28;
        mem[14'd8480] <= 32'hbc8b8403;
        mem[14'd8481] <= 32'hbe48e1a4;
        mem[14'd8482] <= 32'hbe9535fe;
        mem[14'd8483] <= 32'hbea1d49a;
        mem[14'd8484] <= 32'hbe3d25e9;
        mem[14'd8485] <= 32'hbcc74764;
        mem[14'd8486] <= 32'hbb646f84;
        mem[14'd8487] <= 32'hbba0a303;
        mem[14'd8488] <= 32'h3c509ae1;
        mem[14'd8489] <= 32'h3ca0881b;
        mem[14'd8490] <= 32'hbc7f54c7;
        mem[14'd8491] <= 32'hbd9a2de1;
        mem[14'd8492] <= 32'hbe19cab5;
        mem[14'd8493] <= 32'hbe47a83d;
        mem[14'd8494] <= 32'hbe1ce369;
        mem[14'd8495] <= 32'hbe042424;
        mem[14'd8496] <= 32'hbe33c5bb;
        mem[14'd8497] <= 32'hbe8e36a5;
        mem[14'd8498] <= 32'hbe68e5f1;
        mem[14'd8499] <= 32'hbe914e63;
        mem[14'd8500] <= 32'hbe85d218;
        mem[14'd8501] <= 32'hbe30d71c;
        mem[14'd8502] <= 32'hbe305a34;
        mem[14'd8503] <= 32'hbe53c03e;
        mem[14'd8504] <= 32'hbe10c68a;
        mem[14'd8505] <= 32'hbe4c2163;
        mem[14'd8506] <= 32'hbe1db495;
        mem[14'd8507] <= 32'h38565375;
        mem[14'd8508] <= 32'hbceb81b7;
        mem[14'd8509] <= 32'hbe5c1e22;
        mem[14'd8510] <= 32'hbe622467;
        mem[14'd8511] <= 32'hbe4b11d3;
        mem[14'd8512] <= 32'hbda7a754;
        mem[14'd8513] <= 32'hbc8f83c8;
        mem[14'd8514] <= 32'h3b0ebd71;
        mem[14'd8515] <= 32'h3b3cb8c2;
        mem[14'd8516] <= 32'h3ba7631e;
        mem[14'd8517] <= 32'h3bb0a35c;
        mem[14'd8518] <= 32'hbc0a08e5;
        mem[14'd8519] <= 32'hbd8dc081;
        mem[14'd8520] <= 32'hbdefe3d8;
        mem[14'd8521] <= 32'hbdb8371e;
        mem[14'd8522] <= 32'hbe35bbd0;
        mem[14'd8523] <= 32'hbe870c41;
        mem[14'd8524] <= 32'hbe9deb03;
        mem[14'd8525] <= 32'hbed2b097;
        mem[14'd8526] <= 32'hbef814f1;
        mem[14'd8527] <= 32'hbf09d683;
        mem[14'd8528] <= 32'hbf04d304;
        mem[14'd8529] <= 32'hbe6560d3;
        mem[14'd8530] <= 32'hbe8f63d3;
        mem[14'd8531] <= 32'hbe80158a;
        mem[14'd8532] <= 32'hbde2bc27;
        mem[14'd8533] <= 32'hbe224e70;
        mem[14'd8534] <= 32'hbe5240a8;
        mem[14'd8535] <= 32'hbd6399da;
        mem[14'd8536] <= 32'hbddf162b;
        mem[14'd8537] <= 32'hbe7e796b;
        mem[14'd8538] <= 32'hbe2766e4;
        mem[14'd8539] <= 32'hbdb1b959;
        mem[14'd8540] <= 32'h3c29d141;
        mem[14'd8541] <= 32'h3c8b19d8;
        mem[14'd8542] <= 32'hbc3cb0a0;
        mem[14'd8543] <= 32'h3b8b00cb;
        mem[14'd8544] <= 32'h3c0384c7;
        mem[14'd8545] <= 32'h3bb3efc1;
        mem[14'd8546] <= 32'hbbb5053e;
        mem[14'd8547] <= 32'hbdad067b;
        mem[14'd8548] <= 32'hbd94bbe3;
        mem[14'd8549] <= 32'hbda72e54;
        mem[14'd8550] <= 32'hbe055218;
        mem[14'd8551] <= 32'hbe51e112;
        mem[14'd8552] <= 32'hbe5cc59b;
        mem[14'd8553] <= 32'hbe53a947;
        mem[14'd8554] <= 32'hbe7dfabc;
        mem[14'd8555] <= 32'hbeb9425d;
        mem[14'd8556] <= 32'hbea22739;
        mem[14'd8557] <= 32'hbe924397;
        mem[14'd8558] <= 32'hbe9193d0;
        mem[14'd8559] <= 32'hbe76d215;
        mem[14'd8560] <= 32'hbe2cff0d;
        mem[14'd8561] <= 32'hbe8e1e52;
        mem[14'd8562] <= 32'hbe8a78a4;
        mem[14'd8563] <= 32'hbe4c508b;
        mem[14'd8564] <= 32'hbe195094;
        mem[14'd8565] <= 32'hbddc2423;
        mem[14'd8566] <= 32'hbdb198f8;
        mem[14'd8567] <= 32'hbc426fba;
        mem[14'd8568] <= 32'h3d1ad2c8;
        mem[14'd8569] <= 32'hbb7fecc3;
        mem[14'd8570] <= 32'h3bb663a1;
        mem[14'd8571] <= 32'hb9630b48;
        mem[14'd8572] <= 32'h3bc8159f;
        mem[14'd8573] <= 32'hbc4aa747;
        mem[14'd8574] <= 32'h3a55745a;
        mem[14'd8575] <= 32'hbcda8d08;
        mem[14'd8576] <= 32'hbd8195db;
        mem[14'd8577] <= 32'hbe20f47e;
        mem[14'd8578] <= 32'hbe3da0c0;
        mem[14'd8579] <= 32'hbe5cf352;
        mem[14'd8580] <= 32'hbd99878b;
        mem[14'd8581] <= 32'hbdc2b7cb;
        mem[14'd8582] <= 32'hbd2718f1;
        mem[14'd8583] <= 32'hbd29adba;
        mem[14'd8584] <= 32'hbc0a0584;
        mem[14'd8585] <= 32'hbe06122c;
        mem[14'd8586] <= 32'hbd310631;
        mem[14'd8587] <= 32'hbe5cae84;
        mem[14'd8588] <= 32'hbe2f9293;
        mem[14'd8589] <= 32'hbe63908f;
        mem[14'd8590] <= 32'hbe8c4545;
        mem[14'd8591] <= 32'hbeb677cb;
        mem[14'd8592] <= 32'hbdd3e890;
        mem[14'd8593] <= 32'hbd3912a9;
        mem[14'd8594] <= 32'h3d5d6758;
        mem[14'd8595] <= 32'h3da90ac0;
        mem[14'd8596] <= 32'h3d032b25;
        mem[14'd8597] <= 32'hbb2a5c76;
        mem[14'd8598] <= 32'h3bd090d8;
        mem[14'd8599] <= 32'hbbbf3214;
        mem[14'd8600] <= 32'hbbd1456a;
        mem[14'd8601] <= 32'h3bd9417e;
        mem[14'd8602] <= 32'hbbd7c22d;
        mem[14'd8603] <= 32'hbc17cf74;
        mem[14'd8604] <= 32'hbda23d9e;
        mem[14'd8605] <= 32'hbdf5620e;
        mem[14'd8606] <= 32'hbe1ef00c;
        mem[14'd8607] <= 32'hbe21a16e;
        mem[14'd8608] <= 32'h3bdf74f3;
        mem[14'd8609] <= 32'hbe26aef2;
        mem[14'd8610] <= 32'hbd7b038a;
        mem[14'd8611] <= 32'hbdc191ea;
        mem[14'd8612] <= 32'hbdf5dae3;
        mem[14'd8613] <= 32'hbde43c3f;
        mem[14'd8614] <= 32'hbd1e650f;
        mem[14'd8615] <= 32'hbe3086df;
        mem[14'd8616] <= 32'hbe19aacc;
        mem[14'd8617] <= 32'hbe1bb349;
        mem[14'd8618] <= 32'hbe2d6dcc;
        mem[14'd8619] <= 32'hbdeb7dab;
        mem[14'd8620] <= 32'h3cf0711c;
        mem[14'd8621] <= 32'h3e22fce3;
        mem[14'd8622] <= 32'h3e6e7519;
        mem[14'd8623] <= 32'h3e256640;
        mem[14'd8624] <= 32'h3d4fe707;
        mem[14'd8625] <= 32'h3bb15350;
        mem[14'd8626] <= 32'hbc7ca7c9;
        mem[14'd8627] <= 32'hb9c5e587;
        mem[14'd8628] <= 32'hbafa9040;
        mem[14'd8629] <= 32'h3c0c66ed;
        mem[14'd8630] <= 32'hba8a5007;
        mem[14'd8631] <= 32'hbca5af7d;
        mem[14'd8632] <= 32'hbc8af2f5;
        mem[14'd8633] <= 32'h3cc634fe;
        mem[14'd8634] <= 32'h3c9b3e48;
        mem[14'd8635] <= 32'h3db990c0;
        mem[14'd8636] <= 32'h3dc9d60f;
        mem[14'd8637] <= 32'hbdb6b2de;
        mem[14'd8638] <= 32'h3c40599b;
        mem[14'd8639] <= 32'hbdc2a540;
        mem[14'd8640] <= 32'hbe14cad1;
        mem[14'd8641] <= 32'hbe8034c2;
        mem[14'd8642] <= 32'hbe871469;
        mem[14'd8643] <= 32'hbd57aedd;
        mem[14'd8644] <= 32'hbcb2f7c8;
        mem[14'd8645] <= 32'h3d8a6554;
        mem[14'd8646] <= 32'h3d40876b;
        mem[14'd8647] <= 32'h3dfdb766;
        mem[14'd8648] <= 32'h3e912b99;
        mem[14'd8649] <= 32'h3e9dd525;
        mem[14'd8650] <= 32'h3e61acc9;
        mem[14'd8651] <= 32'h3e08774a;
        mem[14'd8652] <= 32'h3c1ff205;
        mem[14'd8653] <= 32'hbc37d9e7;
        mem[14'd8654] <= 32'hbc265ffe;
        mem[14'd8655] <= 32'hbb99838b;
        mem[14'd8656] <= 32'h3caef84b;
        mem[14'd8657] <= 32'h3b83434e;
        mem[14'd8658] <= 32'hbabd5259;
        mem[14'd8659] <= 32'hbc7479aa;
        mem[14'd8660] <= 32'h3bfff323;
        mem[14'd8661] <= 32'h3dffe1a9;
        mem[14'd8662] <= 32'h3e1491fe;
        mem[14'd8663] <= 32'h3e5a5dd3;
        mem[14'd8664] <= 32'h3e789728;
        mem[14'd8665] <= 32'h3e19a242;
        mem[14'd8666] <= 32'h3e5bf1a5;
        mem[14'd8667] <= 32'h3dd5b49f;
        mem[14'd8668] <= 32'h3e2dc4ab;
        mem[14'd8669] <= 32'h3e14b968;
        mem[14'd8670] <= 32'h3e68cbf8;
        mem[14'd8671] <= 32'h3e01d462;
        mem[14'd8672] <= 32'h3e49afdc;
        mem[14'd8673] <= 32'h3e7dd421;
        mem[14'd8674] <= 32'h3ea4ee45;
        mem[14'd8675] <= 32'h3eba2a3b;
        mem[14'd8676] <= 32'h3edef8a5;
        mem[14'd8677] <= 32'h3e9813f4;
        mem[14'd8678] <= 32'h3e0e9930;
        mem[14'd8679] <= 32'h3d24d483;
        mem[14'd8680] <= 32'hbd2c6f7a;
        mem[14'd8681] <= 32'hbc6e751d;
        mem[14'd8682] <= 32'hbc4081d6;
        mem[14'd8683] <= 32'h3c629173;
        mem[14'd8684] <= 32'hbc8dbfbf;
        mem[14'd8685] <= 32'h3bb11c9b;
        mem[14'd8686] <= 32'h3c8e2b98;
        mem[14'd8687] <= 32'hbb8fd5f5;
        mem[14'd8688] <= 32'h3d385039;
        mem[14'd8689] <= 32'h3db15e19;
        mem[14'd8690] <= 32'h3e1ae735;
        mem[14'd8691] <= 32'h3e3b4734;
        mem[14'd8692] <= 32'h3e4b5df8;
        mem[14'd8693] <= 32'h3e9cba89;
        mem[14'd8694] <= 32'h3e9dd61e;
        mem[14'd8695] <= 32'h3ea2bb32;
        mem[14'd8696] <= 32'h3ed04fbe;
        mem[14'd8697] <= 32'h3ec747cd;
        mem[14'd8698] <= 32'h3f01af6f;
        mem[14'd8699] <= 32'h3e9d78cb;
        mem[14'd8700] <= 32'h3e828f3d;
        mem[14'd8701] <= 32'h3e5c6e10;
        mem[14'd8702] <= 32'h3e7a5ebd;
        mem[14'd8703] <= 32'h3e2a4b99;
        mem[14'd8704] <= 32'h3e2e43af;
        mem[14'd8705] <= 32'h3dfd29c3;
        mem[14'd8706] <= 32'h3d008f18;
        mem[14'd8707] <= 32'h3c8c4876;
        mem[14'd8708] <= 32'hbc9ec213;
        mem[14'd8709] <= 32'h3c440b96;
        mem[14'd8710] <= 32'hbbb6e100;
        mem[14'd8711] <= 32'h3c55b761;
        mem[14'd8712] <= 32'hbbb4c9f5;
        mem[14'd8713] <= 32'hbb5271cf;
        mem[14'd8714] <= 32'h3b9c2ccd;
        mem[14'd8715] <= 32'hbb98e098;
        mem[14'd8716] <= 32'hbc24d843;
        mem[14'd8717] <= 32'h3bfe9f19;
        mem[14'd8718] <= 32'hbb4cfa98;
        mem[14'd8719] <= 32'h3c9c6ac9;
        mem[14'd8720] <= 32'h3cb44416;
        mem[14'd8721] <= 32'h3c5cde82;
        mem[14'd8722] <= 32'h3b78e90b;
        mem[14'd8723] <= 32'hbbeb7228;
        mem[14'd8724] <= 32'hba87f46b;
        mem[14'd8725] <= 32'hbd59cf23;
        mem[14'd8726] <= 32'hbc505064;
        mem[14'd8727] <= 32'hbc4e7d53;
        mem[14'd8728] <= 32'hbca71e24;
        mem[14'd8729] <= 32'hbd2c7831;
        mem[14'd8730] <= 32'hbcfd4797;
        mem[14'd8731] <= 32'hbc823a93;
        mem[14'd8732] <= 32'h3bb921b9;
        mem[14'd8733] <= 32'hbc6dd927;
        mem[14'd8734] <= 32'hbc3d0f97;
        mem[14'd8735] <= 32'h3c4eafef;
        mem[14'd8736] <= 32'h3babd512;
        mem[14'd8737] <= 32'hba551f93;
        mem[14'd8738] <= 32'h3b110639;
        mem[14'd8739] <= 32'h3a584e75;
    end

endmodule
