/******************************************************************************
 ** Logisim goes FPGA automatic generated Verilog code                       **
 **                                                                          **
 ** Component : ControllerSignal                                             **
 **                                                                          **
 ******************************************************************************/

`timescale 1ns/1ps
module ControllerSignal( F12,
                         F13,
                         F14,
                         F25,
                         F30,
                         OP2,
                         OP3,
                         OP4,
                         OP5,
                         OP6,
                         ALU_SRC,
                         BEQ,
                         BGE,
                         BLT,
                         BNE,
                         CSRRCI,
                         CSRRSI,
                         FCAL,
                         FLT,
                         FLW,
                         FS0,
                         FS1,
                         FSW,
                         JAL,
                         JALR,
                         LHU,
                         LUI,
                         MemToReg,
                         MemWrite,
                         RegWrite,
                         S_Type,
                         ecall,
                         frd,
                         frs1,
                         frs2,
                         rs1_used,
                         rs2_used);

   /***************************************************************************
    ** Here the inputs are defined                                           **
    ***************************************************************************/
   input  F12;
   input  F13;
   input  F14;
   input  F25;
   input  F30;
   input  OP2;
   input  OP3;
   input  OP4;
   input  OP5;
   input  OP6;

   /***************************************************************************
    ** Here the outputs are defined                                          **
    ***************************************************************************/
   output ALU_SRC;
   output BEQ;
   output BGE;
   output BLT;
   output BNE;
   output CSRRCI;
   output CSRRSI;
   output FCAL;
   output FLT;
   output FLW;
   output FS0;
   output FS1;
   output FSW;
   output JAL;
   output JALR;
   output LHU;
   output LUI;
   output MemToReg;
   output MemWrite;
   output RegWrite;
   output S_Type;
   output ecall;
   output frd;
   output frs1;
   output frs2;
   output rs1_used;
   output rs2_used;

   /***************************************************************************
    ** Here the internal wires are defined                                   **
    ***************************************************************************/
   wire s_LOGISIM_NET_0;
   wire s_LOGISIM_NET_1;
   wire s_LOGISIM_NET_10;
   wire s_LOGISIM_NET_100;
   wire s_LOGISIM_NET_101;
   wire s_LOGISIM_NET_102;
   wire s_LOGISIM_NET_103;
   wire s_LOGISIM_NET_104;
   wire s_LOGISIM_NET_105;
   wire s_LOGISIM_NET_106;
   wire s_LOGISIM_NET_107;
   wire s_LOGISIM_NET_108;
   wire s_LOGISIM_NET_109;
   wire s_LOGISIM_NET_11;
   wire s_LOGISIM_NET_110;
   wire s_LOGISIM_NET_111;
   wire s_LOGISIM_NET_112;
   wire s_LOGISIM_NET_113;
   wire s_LOGISIM_NET_114;
   wire s_LOGISIM_NET_115;
   wire s_LOGISIM_NET_116;
   wire s_LOGISIM_NET_117;
   wire s_LOGISIM_NET_118;
   wire s_LOGISIM_NET_119;
   wire s_LOGISIM_NET_12;
   wire s_LOGISIM_NET_120;
   wire s_LOGISIM_NET_121;
   wire s_LOGISIM_NET_122;
   wire s_LOGISIM_NET_123;
   wire s_LOGISIM_NET_124;
   wire s_LOGISIM_NET_125;
   wire s_LOGISIM_NET_126;
   wire s_LOGISIM_NET_127;
   wire s_LOGISIM_NET_128;
   wire s_LOGISIM_NET_129;
   wire s_LOGISIM_NET_13;
   wire s_LOGISIM_NET_130;
   wire s_LOGISIM_NET_131;
   wire s_LOGISIM_NET_132;
   wire s_LOGISIM_NET_133;
   wire s_LOGISIM_NET_134;
   wire s_LOGISIM_NET_135;
   wire s_LOGISIM_NET_136;
   wire s_LOGISIM_NET_137;
   wire s_LOGISIM_NET_138;
   wire s_LOGISIM_NET_139;
   wire s_LOGISIM_NET_14;
   wire s_LOGISIM_NET_140;
   wire s_LOGISIM_NET_141;
   wire s_LOGISIM_NET_142;
   wire s_LOGISIM_NET_143;
   wire s_LOGISIM_NET_144;
   wire s_LOGISIM_NET_145;
   wire s_LOGISIM_NET_146;
   wire s_LOGISIM_NET_147;
   wire s_LOGISIM_NET_148;
   wire s_LOGISIM_NET_149;
   wire s_LOGISIM_NET_15;
   wire s_LOGISIM_NET_150;
   wire s_LOGISIM_NET_151;
   wire s_LOGISIM_NET_152;
   wire s_LOGISIM_NET_153;
   wire s_LOGISIM_NET_154;
   wire s_LOGISIM_NET_155;
   wire s_LOGISIM_NET_156;
   wire s_LOGISIM_NET_157;
   wire s_LOGISIM_NET_158;
   wire s_LOGISIM_NET_159;
   wire s_LOGISIM_NET_16;
   wire s_LOGISIM_NET_160;
   wire s_LOGISIM_NET_161;
   wire s_LOGISIM_NET_162;
   wire s_LOGISIM_NET_163;
   wire s_LOGISIM_NET_164;
   wire s_LOGISIM_NET_165;
   wire s_LOGISIM_NET_166;
   wire s_LOGISIM_NET_167;
   wire s_LOGISIM_NET_168;
   wire s_LOGISIM_NET_169;
   wire s_LOGISIM_NET_17;
   wire s_LOGISIM_NET_170;
   wire s_LOGISIM_NET_171;
   wire s_LOGISIM_NET_172;
   wire s_LOGISIM_NET_173;
   wire s_LOGISIM_NET_174;
   wire s_LOGISIM_NET_175;
   wire s_LOGISIM_NET_176;
   wire s_LOGISIM_NET_177;
   wire s_LOGISIM_NET_178;
   wire s_LOGISIM_NET_179;
   wire s_LOGISIM_NET_18;
   wire s_LOGISIM_NET_180;
   wire s_LOGISIM_NET_181;
   wire s_LOGISIM_NET_182;
   wire s_LOGISIM_NET_183;
   wire s_LOGISIM_NET_184;
   wire s_LOGISIM_NET_185;
   wire s_LOGISIM_NET_186;
   wire s_LOGISIM_NET_187;
   wire s_LOGISIM_NET_188;
   wire s_LOGISIM_NET_189;
   wire s_LOGISIM_NET_19;
   wire s_LOGISIM_NET_190;
   wire s_LOGISIM_NET_191;
   wire s_LOGISIM_NET_192;
   wire s_LOGISIM_NET_193;
   wire s_LOGISIM_NET_194;
   wire s_LOGISIM_NET_195;
   wire s_LOGISIM_NET_196;
   wire s_LOGISIM_NET_197;
   wire s_LOGISIM_NET_198;
   wire s_LOGISIM_NET_199;
   wire s_LOGISIM_NET_2;
   wire s_LOGISIM_NET_20;
   wire s_LOGISIM_NET_200;
   wire s_LOGISIM_NET_201;
   wire s_LOGISIM_NET_202;
   wire s_LOGISIM_NET_203;
   wire s_LOGISIM_NET_204;
   wire s_LOGISIM_NET_205;
   wire s_LOGISIM_NET_206;
   wire s_LOGISIM_NET_207;
   wire s_LOGISIM_NET_208;
   wire s_LOGISIM_NET_209;
   wire s_LOGISIM_NET_21;
   wire s_LOGISIM_NET_210;
   wire s_LOGISIM_NET_211;
   wire s_LOGISIM_NET_212;
   wire s_LOGISIM_NET_213;
   wire s_LOGISIM_NET_214;
   wire s_LOGISIM_NET_215;
   wire s_LOGISIM_NET_216;
   wire s_LOGISIM_NET_217;
   wire s_LOGISIM_NET_218;
   wire s_LOGISIM_NET_219;
   wire s_LOGISIM_NET_22;
   wire s_LOGISIM_NET_220;
   wire s_LOGISIM_NET_221;
   wire s_LOGISIM_NET_222;
   wire s_LOGISIM_NET_223;
   wire s_LOGISIM_NET_224;
   wire s_LOGISIM_NET_225;
   wire s_LOGISIM_NET_226;
   wire s_LOGISIM_NET_227;
   wire s_LOGISIM_NET_228;
   wire s_LOGISIM_NET_229;
   wire s_LOGISIM_NET_23;
   wire s_LOGISIM_NET_230;
   wire s_LOGISIM_NET_231;
   wire s_LOGISIM_NET_232;
   wire s_LOGISIM_NET_233;
   wire s_LOGISIM_NET_234;
   wire s_LOGISIM_NET_235;
   wire s_LOGISIM_NET_236;
   wire s_LOGISIM_NET_237;
   wire s_LOGISIM_NET_238;
   wire s_LOGISIM_NET_239;
   wire s_LOGISIM_NET_24;
   wire s_LOGISIM_NET_240;
   wire s_LOGISIM_NET_241;
   wire s_LOGISIM_NET_242;
   wire s_LOGISIM_NET_243;
   wire s_LOGISIM_NET_244;
   wire s_LOGISIM_NET_245;
   wire s_LOGISIM_NET_246;
   wire s_LOGISIM_NET_247;
   wire s_LOGISIM_NET_248;
   wire s_LOGISIM_NET_249;
   wire s_LOGISIM_NET_25;
   wire s_LOGISIM_NET_250;
   wire s_LOGISIM_NET_251;
   wire s_LOGISIM_NET_252;
   wire s_LOGISIM_NET_253;
   wire s_LOGISIM_NET_254;
   wire s_LOGISIM_NET_255;
   wire s_LOGISIM_NET_256;
   wire s_LOGISIM_NET_257;
   wire s_LOGISIM_NET_258;
   wire s_LOGISIM_NET_259;
   wire s_LOGISIM_NET_26;
   wire s_LOGISIM_NET_260;
   wire s_LOGISIM_NET_261;
   wire s_LOGISIM_NET_262;
   wire s_LOGISIM_NET_263;
   wire s_LOGISIM_NET_264;
   wire s_LOGISIM_NET_265;
   wire s_LOGISIM_NET_266;
   wire s_LOGISIM_NET_267;
   wire s_LOGISIM_NET_268;
   wire s_LOGISIM_NET_269;
   wire s_LOGISIM_NET_27;
   wire s_LOGISIM_NET_270;
   wire s_LOGISIM_NET_271;
   wire s_LOGISIM_NET_272;
   wire s_LOGISIM_NET_273;
   wire s_LOGISIM_NET_274;
   wire s_LOGISIM_NET_275;
   wire s_LOGISIM_NET_276;
   wire s_LOGISIM_NET_277;
   wire s_LOGISIM_NET_278;
   wire s_LOGISIM_NET_279;
   wire s_LOGISIM_NET_28;
   wire s_LOGISIM_NET_280;
   wire s_LOGISIM_NET_281;
   wire s_LOGISIM_NET_282;
   wire s_LOGISIM_NET_283;
   wire s_LOGISIM_NET_284;
   wire s_LOGISIM_NET_285;
   wire s_LOGISIM_NET_286;
   wire s_LOGISIM_NET_287;
   wire s_LOGISIM_NET_288;
   wire s_LOGISIM_NET_289;
   wire s_LOGISIM_NET_29;
   wire s_LOGISIM_NET_290;
   wire s_LOGISIM_NET_291;
   wire s_LOGISIM_NET_292;
   wire s_LOGISIM_NET_293;
   wire s_LOGISIM_NET_294;
   wire s_LOGISIM_NET_295;
   wire s_LOGISIM_NET_296;
   wire s_LOGISIM_NET_297;
   wire s_LOGISIM_NET_298;
   wire s_LOGISIM_NET_299;
   wire s_LOGISIM_NET_3;
   wire s_LOGISIM_NET_30;
   wire s_LOGISIM_NET_300;
   wire s_LOGISIM_NET_301;
   wire s_LOGISIM_NET_302;
   wire s_LOGISIM_NET_303;
   wire s_LOGISIM_NET_304;
   wire s_LOGISIM_NET_305;
   wire s_LOGISIM_NET_306;
   wire s_LOGISIM_NET_307;
   wire s_LOGISIM_NET_308;
   wire s_LOGISIM_NET_309;
   wire s_LOGISIM_NET_31;
   wire s_LOGISIM_NET_310;
   wire s_LOGISIM_NET_311;
   wire s_LOGISIM_NET_312;
   wire s_LOGISIM_NET_313;
   wire s_LOGISIM_NET_314;
   wire s_LOGISIM_NET_315;
   wire s_LOGISIM_NET_316;
   wire s_LOGISIM_NET_317;
   wire s_LOGISIM_NET_318;
   wire s_LOGISIM_NET_319;
   wire s_LOGISIM_NET_32;
   wire s_LOGISIM_NET_320;
   wire s_LOGISIM_NET_321;
   wire s_LOGISIM_NET_322;
   wire s_LOGISIM_NET_323;
   wire s_LOGISIM_NET_324;
   wire s_LOGISIM_NET_325;
   wire s_LOGISIM_NET_326;
   wire s_LOGISIM_NET_327;
   wire s_LOGISIM_NET_328;
   wire s_LOGISIM_NET_329;
   wire s_LOGISIM_NET_33;
   wire s_LOGISIM_NET_330;
   wire s_LOGISIM_NET_331;
   wire s_LOGISIM_NET_332;
   wire s_LOGISIM_NET_333;
   wire s_LOGISIM_NET_334;
   wire s_LOGISIM_NET_335;
   wire s_LOGISIM_NET_336;
   wire s_LOGISIM_NET_337;
   wire s_LOGISIM_NET_338;
   wire s_LOGISIM_NET_339;
   wire s_LOGISIM_NET_34;
   wire s_LOGISIM_NET_340;
   wire s_LOGISIM_NET_341;
   wire s_LOGISIM_NET_342;
   wire s_LOGISIM_NET_343;
   wire s_LOGISIM_NET_344;
   wire s_LOGISIM_NET_345;
   wire s_LOGISIM_NET_346;
   wire s_LOGISIM_NET_347;
   wire s_LOGISIM_NET_348;
   wire s_LOGISIM_NET_349;
   wire s_LOGISIM_NET_35;
   wire s_LOGISIM_NET_350;
   wire s_LOGISIM_NET_351;
   wire s_LOGISIM_NET_352;
   wire s_LOGISIM_NET_353;
   wire s_LOGISIM_NET_354;
   wire s_LOGISIM_NET_355;
   wire s_LOGISIM_NET_356;
   wire s_LOGISIM_NET_357;
   wire s_LOGISIM_NET_358;
   wire s_LOGISIM_NET_359;
   wire s_LOGISIM_NET_36;
   wire s_LOGISIM_NET_360;
   wire s_LOGISIM_NET_361;
   wire s_LOGISIM_NET_362;
   wire s_LOGISIM_NET_363;
   wire s_LOGISIM_NET_364;
   wire s_LOGISIM_NET_365;
   wire s_LOGISIM_NET_366;
   wire s_LOGISIM_NET_367;
   wire s_LOGISIM_NET_368;
   wire s_LOGISIM_NET_369;
   wire s_LOGISIM_NET_37;
   wire s_LOGISIM_NET_370;
   wire s_LOGISIM_NET_371;
   wire s_LOGISIM_NET_372;
   wire s_LOGISIM_NET_373;
   wire s_LOGISIM_NET_374;
   wire s_LOGISIM_NET_375;
   wire s_LOGISIM_NET_376;
   wire s_LOGISIM_NET_377;
   wire s_LOGISIM_NET_378;
   wire s_LOGISIM_NET_379;
   wire s_LOGISIM_NET_38;
   wire s_LOGISIM_NET_380;
   wire s_LOGISIM_NET_381;
   wire s_LOGISIM_NET_382;
   wire s_LOGISIM_NET_383;
   wire s_LOGISIM_NET_384;
   wire s_LOGISIM_NET_385;
   wire s_LOGISIM_NET_386;
   wire s_LOGISIM_NET_387;
   wire s_LOGISIM_NET_388;
   wire s_LOGISIM_NET_389;
   wire s_LOGISIM_NET_39;
   wire s_LOGISIM_NET_390;
   wire s_LOGISIM_NET_391;
   wire s_LOGISIM_NET_392;
   wire s_LOGISIM_NET_393;
   wire s_LOGISIM_NET_394;
   wire s_LOGISIM_NET_395;
   wire s_LOGISIM_NET_396;
   wire s_LOGISIM_NET_397;
   wire s_LOGISIM_NET_398;
   wire s_LOGISIM_NET_399;
   wire s_LOGISIM_NET_4;
   wire s_LOGISIM_NET_40;
   wire s_LOGISIM_NET_400;
   wire s_LOGISIM_NET_401;
   wire s_LOGISIM_NET_402;
   wire s_LOGISIM_NET_403;
   wire s_LOGISIM_NET_404;
   wire s_LOGISIM_NET_405;
   wire s_LOGISIM_NET_406;
   wire s_LOGISIM_NET_407;
   wire s_LOGISIM_NET_408;
   wire s_LOGISIM_NET_409;
   wire s_LOGISIM_NET_41;
   wire s_LOGISIM_NET_410;
   wire s_LOGISIM_NET_411;
   wire s_LOGISIM_NET_412;
   wire s_LOGISIM_NET_413;
   wire s_LOGISIM_NET_414;
   wire s_LOGISIM_NET_415;
   wire s_LOGISIM_NET_416;
   wire s_LOGISIM_NET_417;
   wire s_LOGISIM_NET_418;
   wire s_LOGISIM_NET_419;
   wire s_LOGISIM_NET_42;
   wire s_LOGISIM_NET_420;
   wire s_LOGISIM_NET_421;
   wire s_LOGISIM_NET_422;
   wire s_LOGISIM_NET_423;
   wire s_LOGISIM_NET_424;
   wire s_LOGISIM_NET_425;
   wire s_LOGISIM_NET_426;
   wire s_LOGISIM_NET_427;
   wire s_LOGISIM_NET_428;
   wire s_LOGISIM_NET_429;
   wire s_LOGISIM_NET_43;
   wire s_LOGISIM_NET_430;
   wire s_LOGISIM_NET_431;
   wire s_LOGISIM_NET_432;
   wire s_LOGISIM_NET_433;
   wire s_LOGISIM_NET_434;
   wire s_LOGISIM_NET_435;
   wire s_LOGISIM_NET_436;
   wire s_LOGISIM_NET_437;
   wire s_LOGISIM_NET_438;
   wire s_LOGISIM_NET_439;
   wire s_LOGISIM_NET_44;
   wire s_LOGISIM_NET_440;
   wire s_LOGISIM_NET_441;
   wire s_LOGISIM_NET_442;
   wire s_LOGISIM_NET_443;
   wire s_LOGISIM_NET_444;
   wire s_LOGISIM_NET_445;
   wire s_LOGISIM_NET_446;
   wire s_LOGISIM_NET_447;
   wire s_LOGISIM_NET_448;
   wire s_LOGISIM_NET_449;
   wire s_LOGISIM_NET_45;
   wire s_LOGISIM_NET_450;
   wire s_LOGISIM_NET_451;
   wire s_LOGISIM_NET_452;
   wire s_LOGISIM_NET_453;
   wire s_LOGISIM_NET_454;
   wire s_LOGISIM_NET_455;
   wire s_LOGISIM_NET_456;
   wire s_LOGISIM_NET_457;
   wire s_LOGISIM_NET_458;
   wire s_LOGISIM_NET_459;
   wire s_LOGISIM_NET_46;
   wire s_LOGISIM_NET_460;
   wire s_LOGISIM_NET_461;
   wire s_LOGISIM_NET_462;
   wire s_LOGISIM_NET_463;
   wire s_LOGISIM_NET_464;
   wire s_LOGISIM_NET_465;
   wire s_LOGISIM_NET_466;
   wire s_LOGISIM_NET_467;
   wire s_LOGISIM_NET_468;
   wire s_LOGISIM_NET_469;
   wire s_LOGISIM_NET_47;
   wire s_LOGISIM_NET_470;
   wire s_LOGISIM_NET_471;
   wire s_LOGISIM_NET_472;
   wire s_LOGISIM_NET_473;
   wire s_LOGISIM_NET_474;
   wire s_LOGISIM_NET_475;
   wire s_LOGISIM_NET_476;
   wire s_LOGISIM_NET_477;
   wire s_LOGISIM_NET_478;
   wire s_LOGISIM_NET_479;
   wire s_LOGISIM_NET_48;
   wire s_LOGISIM_NET_480;
   wire s_LOGISIM_NET_481;
   wire s_LOGISIM_NET_482;
   wire s_LOGISIM_NET_483;
   wire s_LOGISIM_NET_484;
   wire s_LOGISIM_NET_485;
   wire s_LOGISIM_NET_486;
   wire s_LOGISIM_NET_487;
   wire s_LOGISIM_NET_488;
   wire s_LOGISIM_NET_489;
   wire s_LOGISIM_NET_49;
   wire s_LOGISIM_NET_490;
   wire s_LOGISIM_NET_491;
   wire s_LOGISIM_NET_492;
   wire s_LOGISIM_NET_493;
   wire s_LOGISIM_NET_494;
   wire s_LOGISIM_NET_495;
   wire s_LOGISIM_NET_496;
   wire s_LOGISIM_NET_497;
   wire s_LOGISIM_NET_498;
   wire s_LOGISIM_NET_499;
   wire s_LOGISIM_NET_5;
   wire s_LOGISIM_NET_50;
   wire s_LOGISIM_NET_500;
   wire s_LOGISIM_NET_501;
   wire s_LOGISIM_NET_502;
   wire s_LOGISIM_NET_503;
   wire s_LOGISIM_NET_504;
   wire s_LOGISIM_NET_505;
   wire s_LOGISIM_NET_506;
   wire s_LOGISIM_NET_507;
   wire s_LOGISIM_NET_508;
   wire s_LOGISIM_NET_509;
   wire s_LOGISIM_NET_51;
   wire s_LOGISIM_NET_510;
   wire s_LOGISIM_NET_511;
   wire s_LOGISIM_NET_512;
   wire s_LOGISIM_NET_513;
   wire s_LOGISIM_NET_514;
   wire s_LOGISIM_NET_515;
   wire s_LOGISIM_NET_516;
   wire s_LOGISIM_NET_517;
   wire s_LOGISIM_NET_518;
   wire s_LOGISIM_NET_519;
   wire s_LOGISIM_NET_52;
   wire s_LOGISIM_NET_520;
   wire s_LOGISIM_NET_521;
   wire s_LOGISIM_NET_522;
   wire s_LOGISIM_NET_523;
   wire s_LOGISIM_NET_524;
   wire s_LOGISIM_NET_525;
   wire s_LOGISIM_NET_526;
   wire s_LOGISIM_NET_527;
   wire s_LOGISIM_NET_528;
   wire s_LOGISIM_NET_529;
   wire s_LOGISIM_NET_53;
   wire s_LOGISIM_NET_530;
   wire s_LOGISIM_NET_531;
   wire s_LOGISIM_NET_532;
   wire s_LOGISIM_NET_533;
   wire s_LOGISIM_NET_534;
   wire s_LOGISIM_NET_535;
   wire s_LOGISIM_NET_536;
   wire s_LOGISIM_NET_537;
   wire s_LOGISIM_NET_538;
   wire s_LOGISIM_NET_539;
   wire s_LOGISIM_NET_54;
   wire s_LOGISIM_NET_540;
   wire s_LOGISIM_NET_541;
   wire s_LOGISIM_NET_542;
   wire s_LOGISIM_NET_543;
   wire s_LOGISIM_NET_544;
   wire s_LOGISIM_NET_545;
   wire s_LOGISIM_NET_546;
   wire s_LOGISIM_NET_547;
   wire s_LOGISIM_NET_548;
   wire s_LOGISIM_NET_549;
   wire s_LOGISIM_NET_55;
   wire s_LOGISIM_NET_550;
   wire s_LOGISIM_NET_551;
   wire s_LOGISIM_NET_552;
   wire s_LOGISIM_NET_553;
   wire s_LOGISIM_NET_554;
   wire s_LOGISIM_NET_555;
   wire s_LOGISIM_NET_556;
   wire s_LOGISIM_NET_557;
   wire s_LOGISIM_NET_558;
   wire s_LOGISIM_NET_559;
   wire s_LOGISIM_NET_56;
   wire s_LOGISIM_NET_560;
   wire s_LOGISIM_NET_561;
   wire s_LOGISIM_NET_562;
   wire s_LOGISIM_NET_563;
   wire s_LOGISIM_NET_564;
   wire s_LOGISIM_NET_565;
   wire s_LOGISIM_NET_566;
   wire s_LOGISIM_NET_567;
   wire s_LOGISIM_NET_568;
   wire s_LOGISIM_NET_569;
   wire s_LOGISIM_NET_57;
   wire s_LOGISIM_NET_570;
   wire s_LOGISIM_NET_571;
   wire s_LOGISIM_NET_572;
   wire s_LOGISIM_NET_573;
   wire s_LOGISIM_NET_574;
   wire s_LOGISIM_NET_575;
   wire s_LOGISIM_NET_576;
   wire s_LOGISIM_NET_577;
   wire s_LOGISIM_NET_578;
   wire s_LOGISIM_NET_579;
   wire s_LOGISIM_NET_58;
   wire s_LOGISIM_NET_580;
   wire s_LOGISIM_NET_581;
   wire s_LOGISIM_NET_582;
   wire s_LOGISIM_NET_583;
   wire s_LOGISIM_NET_584;
   wire s_LOGISIM_NET_585;
   wire s_LOGISIM_NET_586;
   wire s_LOGISIM_NET_587;
   wire s_LOGISIM_NET_588;
   wire s_LOGISIM_NET_589;
   wire s_LOGISIM_NET_59;
   wire s_LOGISIM_NET_590;
   wire s_LOGISIM_NET_591;
   wire s_LOGISIM_NET_592;
   wire s_LOGISIM_NET_593;
   wire s_LOGISIM_NET_594;
   wire s_LOGISIM_NET_595;
   wire s_LOGISIM_NET_596;
   wire s_LOGISIM_NET_597;
   wire s_LOGISIM_NET_598;
   wire s_LOGISIM_NET_599;
   wire s_LOGISIM_NET_6;
   wire s_LOGISIM_NET_60;
   wire s_LOGISIM_NET_600;
   wire s_LOGISIM_NET_601;
   wire s_LOGISIM_NET_602;
   wire s_LOGISIM_NET_603;
   wire s_LOGISIM_NET_604;
   wire s_LOGISIM_NET_605;
   wire s_LOGISIM_NET_606;
   wire s_LOGISIM_NET_607;
   wire s_LOGISIM_NET_608;
   wire s_LOGISIM_NET_609;
   wire s_LOGISIM_NET_61;
   wire s_LOGISIM_NET_610;
   wire s_LOGISIM_NET_611;
   wire s_LOGISIM_NET_612;
   wire s_LOGISIM_NET_613;
   wire s_LOGISIM_NET_614;
   wire s_LOGISIM_NET_615;
   wire s_LOGISIM_NET_616;
   wire s_LOGISIM_NET_617;
   wire s_LOGISIM_NET_618;
   wire s_LOGISIM_NET_619;
   wire s_LOGISIM_NET_62;
   wire s_LOGISIM_NET_620;
   wire s_LOGISIM_NET_621;
   wire s_LOGISIM_NET_622;
   wire s_LOGISIM_NET_623;
   wire s_LOGISIM_NET_624;
   wire s_LOGISIM_NET_625;
   wire s_LOGISIM_NET_626;
   wire s_LOGISIM_NET_627;
   wire s_LOGISIM_NET_628;
   wire s_LOGISIM_NET_629;
   wire s_LOGISIM_NET_63;
   wire s_LOGISIM_NET_630;
   wire s_LOGISIM_NET_631;
   wire s_LOGISIM_NET_632;
   wire s_LOGISIM_NET_633;
   wire s_LOGISIM_NET_634;
   wire s_LOGISIM_NET_635;
   wire s_LOGISIM_NET_636;
   wire s_LOGISIM_NET_637;
   wire s_LOGISIM_NET_638;
   wire s_LOGISIM_NET_639;
   wire s_LOGISIM_NET_64;
   wire s_LOGISIM_NET_640;
   wire s_LOGISIM_NET_641;
   wire s_LOGISIM_NET_642;
   wire s_LOGISIM_NET_643;
   wire s_LOGISIM_NET_644;
   wire s_LOGISIM_NET_645;
   wire s_LOGISIM_NET_646;
   wire s_LOGISIM_NET_647;
   wire s_LOGISIM_NET_648;
   wire s_LOGISIM_NET_649;
   wire s_LOGISIM_NET_65;
   wire s_LOGISIM_NET_650;
   wire s_LOGISIM_NET_651;
   wire s_LOGISIM_NET_652;
   wire s_LOGISIM_NET_653;
   wire s_LOGISIM_NET_654;
   wire s_LOGISIM_NET_655;
   wire s_LOGISIM_NET_656;
   wire s_LOGISIM_NET_657;
   wire s_LOGISIM_NET_658;
   wire s_LOGISIM_NET_659;
   wire s_LOGISIM_NET_66;
   wire s_LOGISIM_NET_660;
   wire s_LOGISIM_NET_661;
   wire s_LOGISIM_NET_662;
   wire s_LOGISIM_NET_663;
   wire s_LOGISIM_NET_664;
   wire s_LOGISIM_NET_665;
   wire s_LOGISIM_NET_666;
   wire s_LOGISIM_NET_667;
   wire s_LOGISIM_NET_668;
   wire s_LOGISIM_NET_669;
   wire s_LOGISIM_NET_67;
   wire s_LOGISIM_NET_670;
   wire s_LOGISIM_NET_671;
   wire s_LOGISIM_NET_672;
   wire s_LOGISIM_NET_673;
   wire s_LOGISIM_NET_674;
   wire s_LOGISIM_NET_675;
   wire s_LOGISIM_NET_676;
   wire s_LOGISIM_NET_677;
   wire s_LOGISIM_NET_678;
   wire s_LOGISIM_NET_679;
   wire s_LOGISIM_NET_68;
   wire s_LOGISIM_NET_680;
   wire s_LOGISIM_NET_681;
   wire s_LOGISIM_NET_682;
   wire s_LOGISIM_NET_683;
   wire s_LOGISIM_NET_684;
   wire s_LOGISIM_NET_685;
   wire s_LOGISIM_NET_686;
   wire s_LOGISIM_NET_687;
   wire s_LOGISIM_NET_688;
   wire s_LOGISIM_NET_689;
   wire s_LOGISIM_NET_69;
   wire s_LOGISIM_NET_690;
   wire s_LOGISIM_NET_691;
   wire s_LOGISIM_NET_692;
   wire s_LOGISIM_NET_693;
   wire s_LOGISIM_NET_694;
   wire s_LOGISIM_NET_695;
   wire s_LOGISIM_NET_696;
   wire s_LOGISIM_NET_697;
   wire s_LOGISIM_NET_698;
   wire s_LOGISIM_NET_699;
   wire s_LOGISIM_NET_7;
   wire s_LOGISIM_NET_70;
   wire s_LOGISIM_NET_700;
   wire s_LOGISIM_NET_701;
   wire s_LOGISIM_NET_702;
   wire s_LOGISIM_NET_703;
   wire s_LOGISIM_NET_704;
   wire s_LOGISIM_NET_705;
   wire s_LOGISIM_NET_706;
   wire s_LOGISIM_NET_707;
   wire s_LOGISIM_NET_708;
   wire s_LOGISIM_NET_709;
   wire s_LOGISIM_NET_71;
   wire s_LOGISIM_NET_710;
   wire s_LOGISIM_NET_711;
   wire s_LOGISIM_NET_712;
   wire s_LOGISIM_NET_713;
   wire s_LOGISIM_NET_714;
   wire s_LOGISIM_NET_715;
   wire s_LOGISIM_NET_716;
   wire s_LOGISIM_NET_717;
   wire s_LOGISIM_NET_718;
   wire s_LOGISIM_NET_719;
   wire s_LOGISIM_NET_72;
   wire s_LOGISIM_NET_720;
   wire s_LOGISIM_NET_721;
   wire s_LOGISIM_NET_722;
   wire s_LOGISIM_NET_723;
   wire s_LOGISIM_NET_724;
   wire s_LOGISIM_NET_725;
   wire s_LOGISIM_NET_726;
   wire s_LOGISIM_NET_727;
   wire s_LOGISIM_NET_728;
   wire s_LOGISIM_NET_729;
   wire s_LOGISIM_NET_73;
   wire s_LOGISIM_NET_730;
   wire s_LOGISIM_NET_731;
   wire s_LOGISIM_NET_732;
   wire s_LOGISIM_NET_733;
   wire s_LOGISIM_NET_734;
   wire s_LOGISIM_NET_735;
   wire s_LOGISIM_NET_736;
   wire s_LOGISIM_NET_737;
   wire s_LOGISIM_NET_738;
   wire s_LOGISIM_NET_739;
   wire s_LOGISIM_NET_74;
   wire s_LOGISIM_NET_740;
   wire s_LOGISIM_NET_741;
   wire s_LOGISIM_NET_742;
   wire s_LOGISIM_NET_743;
   wire s_LOGISIM_NET_744;
   wire s_LOGISIM_NET_745;
   wire s_LOGISIM_NET_746;
   wire s_LOGISIM_NET_747;
   wire s_LOGISIM_NET_748;
   wire s_LOGISIM_NET_749;
   wire s_LOGISIM_NET_75;
   wire s_LOGISIM_NET_750;
   wire s_LOGISIM_NET_751;
   wire s_LOGISIM_NET_752;
   wire s_LOGISIM_NET_753;
   wire s_LOGISIM_NET_754;
   wire s_LOGISIM_NET_755;
   wire s_LOGISIM_NET_756;
   wire s_LOGISIM_NET_757;
   wire s_LOGISIM_NET_758;
   wire s_LOGISIM_NET_759;
   wire s_LOGISIM_NET_76;
   wire s_LOGISIM_NET_760;
   wire s_LOGISIM_NET_761;
   wire s_LOGISIM_NET_762;
   wire s_LOGISIM_NET_763;
   wire s_LOGISIM_NET_764;
   wire s_LOGISIM_NET_765;
   wire s_LOGISIM_NET_766;
   wire s_LOGISIM_NET_767;
   wire s_LOGISIM_NET_768;
   wire s_LOGISIM_NET_769;
   wire s_LOGISIM_NET_77;
   wire s_LOGISIM_NET_770;
   wire s_LOGISIM_NET_771;
   wire s_LOGISIM_NET_772;
   wire s_LOGISIM_NET_773;
   wire s_LOGISIM_NET_774;
   wire s_LOGISIM_NET_775;
   wire s_LOGISIM_NET_776;
   wire s_LOGISIM_NET_777;
   wire s_LOGISIM_NET_778;
   wire s_LOGISIM_NET_779;
   wire s_LOGISIM_NET_78;
   wire s_LOGISIM_NET_780;
   wire s_LOGISIM_NET_781;
   wire s_LOGISIM_NET_782;
   wire s_LOGISIM_NET_783;
   wire s_LOGISIM_NET_784;
   wire s_LOGISIM_NET_785;
   wire s_LOGISIM_NET_786;
   wire s_LOGISIM_NET_787;
   wire s_LOGISIM_NET_788;
   wire s_LOGISIM_NET_789;
   wire s_LOGISIM_NET_79;
   wire s_LOGISIM_NET_790;
   wire s_LOGISIM_NET_791;
   wire s_LOGISIM_NET_792;
   wire s_LOGISIM_NET_793;
   wire s_LOGISIM_NET_794;
   wire s_LOGISIM_NET_795;
   wire s_LOGISIM_NET_796;
   wire s_LOGISIM_NET_797;
   wire s_LOGISIM_NET_798;
   wire s_LOGISIM_NET_799;
   wire s_LOGISIM_NET_8;
   wire s_LOGISIM_NET_80;
   wire s_LOGISIM_NET_800;
   wire s_LOGISIM_NET_801;
   wire s_LOGISIM_NET_802;
   wire s_LOGISIM_NET_803;
   wire s_LOGISIM_NET_804;
   wire s_LOGISIM_NET_81;
   wire s_LOGISIM_NET_82;
   wire s_LOGISIM_NET_83;
   wire s_LOGISIM_NET_84;
   wire s_LOGISIM_NET_85;
   wire s_LOGISIM_NET_86;
   wire s_LOGISIM_NET_87;
   wire s_LOGISIM_NET_88;
   wire s_LOGISIM_NET_89;
   wire s_LOGISIM_NET_9;
   wire s_LOGISIM_NET_90;
   wire s_LOGISIM_NET_91;
   wire s_LOGISIM_NET_92;
   wire s_LOGISIM_NET_93;
   wire s_LOGISIM_NET_94;
   wire s_LOGISIM_NET_95;
   wire s_LOGISIM_NET_96;
   wire s_LOGISIM_NET_97;
   wire s_LOGISIM_NET_98;
   wire s_LOGISIM_NET_99;


   /***************************************************************************
    ** Here all input connections are defined                                **
    ***************************************************************************/
   assign s_LOGISIM_NET_17                   = OP2;
   assign s_LOGISIM_NET_7                    = F14;
   assign s_LOGISIM_NET_21                   = OP5;
   assign s_LOGISIM_NET_20                   = F30;
   assign s_LOGISIM_NET_8                    = F12;
   assign s_LOGISIM_NET_54                   = OP6;
   assign s_LOGISIM_NET_10                   = OP3;
   assign s_LOGISIM_NET_3                    = OP4;
   assign s_LOGISIM_NET_1                    = F25;
   assign s_LOGISIM_NET_9                    = F13;

   /***************************************************************************
    ** Here all output connections are defined                               **
    ***************************************************************************/
   assign FLW                                = s_LOGISIM_NET_548;
   assign MemWrite                           = s_LOGISIM_NET_670;
   assign BGE                                = s_LOGISIM_NET_730;
   assign frd                                = s_LOGISIM_NET_766;
   assign JALR                               = s_LOGISIM_NET_734;
   assign FLT                                = s_LOGISIM_NET_397;
   assign frs2                               = s_LOGISIM_NET_736;
   assign FCAL                               = s_LOGISIM_NET_728;
   assign rs1_used                           = s_LOGISIM_NET_15;
   assign LUI                                = s_LOGISIM_NET_190;
   assign FS1                                = s_LOGISIM_NET_733;
   assign LHU                                = s_LOGISIM_NET_791;
   assign ALU_SRC                            = s_LOGISIM_NET_226;
   assign CSRRCI                             = s_LOGISIM_NET_723;
   assign BNE                                = s_LOGISIM_NET_780;
   assign FS0                                = s_LOGISIM_NET_787;
   assign RegWrite                           = s_LOGISIM_NET_68;
   assign BLT                                = s_LOGISIM_NET_219;
   assign MemToReg                           = s_LOGISIM_NET_796;
   assign JAL                                = s_LOGISIM_NET_769;
   assign CSRRSI                             = s_LOGISIM_NET_175;
   assign frs1                               = s_LOGISIM_NET_778;
   assign S_Type                             = s_LOGISIM_NET_324;
   assign FSW                                = s_LOGISIM_NET_740;
   assign rs2_used                           = s_LOGISIM_NET_795;
   assign BEQ                                = s_LOGISIM_NET_192;
   assign ecall                              = s_LOGISIM_NET_804;

   /***************************************************************************
    ** Here all normal components are defined                                **
    ***************************************************************************/
   NOT_GATE      GATE_1 (.Input_1(s_LOGISIM_NET_7),
                         .Result(s_LOGISIM_NET_630));

   NOT_GATE      GATE_2 (.Input_1(s_LOGISIM_NET_54),
                         .Result(s_LOGISIM_NET_557));

   NOT_GATE      GATE_3 (.Input_1(s_LOGISIM_NET_1),
                         .Result(s_LOGISIM_NET_452));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_4 (.Input_1(s_LOGISIM_NET_272),
              .Input_2(s_LOGISIM_NET_9),
              .Input_3(s_LOGISIM_NET_198),
              .Input_4(s_LOGISIM_NET_714),
              .Input_5(s_LOGISIM_NET_63),
              .Input_6(s_LOGISIM_NET_207),
              .Input_7(s_LOGISIM_NET_534),
              .Input_8(s_LOGISIM_NET_17),
              .Result(s_LOGISIM_NET_548));

   NOT_GATE      GATE_5 (.Input_1(s_LOGISIM_NET_1),
                         .Result(s_LOGISIM_NET_732));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_6 (.Input_1(s_LOGISIM_NET_265),
              .Input_10(s_LOGISIM_NET_782),
              .Input_2(s_LOGISIM_NET_164),
              .Input_3(s_LOGISIM_NET_420),
              .Input_4(s_LOGISIM_NET_229),
              .Input_5(s_LOGISIM_NET_8),
              .Input_6(s_LOGISIM_NET_54),
              .Input_7(s_LOGISIM_NET_167),
              .Input_8(s_LOGISIM_NET_3),
              .Input_9(s_LOGISIM_NET_698),
              .Result(s_LOGISIM_NET_421));

   NOT_GATE      GATE_7 (.Input_1(s_LOGISIM_NET_3),
                         .Result(s_LOGISIM_NET_560));

   NOT_GATE      GATE_8 (.Input_1(s_LOGISIM_NET_17),
                         .Result(s_LOGISIM_NET_520));

   NOT_GATE      GATE_9 (.Input_1(s_LOGISIM_NET_21),
                         .Result(s_LOGISIM_NET_158));

   NOT_GATE      GATE_10 (.Input_1(s_LOGISIM_NET_8),
                          .Result(s_LOGISIM_NET_77));

   NOT_GATE      GATE_11 (.Input_1(s_LOGISIM_NET_54),
                          .Result(s_LOGISIM_NET_186));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_12 (.Input_1(s_LOGISIM_NET_7),
               .Input_2(s_LOGISIM_NET_612),
               .Input_3(s_LOGISIM_NET_537),
               .Input_4(s_LOGISIM_NET_54),
               .Input_5(s_LOGISIM_NET_21),
               .Input_6(s_LOGISIM_NET_143),
               .Input_7(s_LOGISIM_NET_400),
               .Input_8(s_LOGISIM_NET_108),
               .Result(s_LOGISIM_NET_507));

   NOT_GATE      GATE_13 (.Input_1(s_LOGISIM_NET_54),
                          .Result(s_LOGISIM_NET_297));

   NOT_GATE      GATE_14 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_441));

   NOT_GATE      GATE_15 (.Input_1(s_LOGISIM_NET_9),
                          .Result(s_LOGISIM_NET_125));

   NOT_GATE      GATE_16 (.Input_1(s_LOGISIM_NET_8),
                          .Result(s_LOGISIM_NET_268));

   NOT_GATE      GATE_17 (.Input_1(s_LOGISIM_NET_8),
                          .Result(s_LOGISIM_NET_352));

   NOT_GATE      GATE_18 (.Input_1(s_LOGISIM_NET_17),
                          .Result(s_LOGISIM_NET_144));

   NOT_GATE      GATE_19 (.Input_1(s_LOGISIM_NET_17),
                          .Result(s_LOGISIM_NET_600));

   NOT_GATE      GATE_20 (.Input_1(s_LOGISIM_NET_21),
                          .Result(s_LOGISIM_NET_748));

   NOT_GATE      GATE_21 (.Input_1(s_LOGISIM_NET_10),
                          .Result(s_LOGISIM_NET_602));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_22 (.Input_1(s_LOGISIM_NET_438),
               .Input_2(s_LOGISIM_NET_320),
               .Input_3(s_LOGISIM_NET_149),
               .Input_4(s_LOGISIM_NET_54),
               .Input_5(s_LOGISIM_NET_21),
               .Input_6(s_LOGISIM_NET_442),
               .Input_7(s_LOGISIM_NET_662),
               .Input_8(s_LOGISIM_NET_205),
               .Result(s_LOGISIM_NET_178));

   NOT_GATE      GATE_23 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_172));

   NOT_GATE      GATE_24 (.Input_1(s_LOGISIM_NET_10),
                          .Result(s_LOGISIM_NET_538));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_25 (.Input_1(s_LOGISIM_NET_7),
               .Input_2(s_LOGISIM_NET_9),
               .Input_3(s_LOGISIM_NET_668),
               .Input_4(s_LOGISIM_NET_453),
               .Input_5(s_LOGISIM_NET_368),
               .Input_6(s_LOGISIM_NET_3),
               .Input_7(s_LOGISIM_NET_11),
               .Input_8(s_LOGISIM_NET_437),
               .Result(s_LOGISIM_NET_422));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_26 (.Input_1(s_LOGISIM_NET_764),
               .Input_2(s_LOGISIM_NET_9),
               .Input_3(s_LOGISIM_NET_644),
               .Input_4(s_LOGISIM_NET_417),
               .Input_5(s_LOGISIM_NET_323),
               .Input_6(s_LOGISIM_NET_3),
               .Input_7(s_LOGISIM_NET_201),
               .Input_8(s_LOGISIM_NET_410),
               .Result(s_LOGISIM_NET_148));

   NOT_GATE      GATE_27 (.Input_1(s_LOGISIM_NET_8),
                          .Result(s_LOGISIM_NET_402));

   NOT_GATE      GATE_28 (.Input_1(s_LOGISIM_NET_8),
                          .Result(s_LOGISIM_NET_328));

   NOT_GATE      GATE_29 (.Input_1(s_LOGISIM_NET_20),
                          .Result(s_LOGISIM_NET_231));

   NOT_GATE      GATE_30 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_76));

   NOT_GATE      GATE_31 (.Input_1(s_LOGISIM_NET_54),
                          .Result(s_LOGISIM_NET_711));

   NOT_GATE      GATE_32 (.Input_1(s_LOGISIM_NET_10),
                          .Result(s_LOGISIM_NET_115));

   NOT_GATE      GATE_33 (.Input_1(s_LOGISIM_NET_10),
                          .Result(s_LOGISIM_NET_136));

   NOT_GATE      GATE_34 (.Input_1(s_LOGISIM_NET_17),
                          .Result(s_LOGISIM_NET_549));

   NOT_GATE      GATE_35 (.Input_1(s_LOGISIM_NET_20),
                          .Result(s_LOGISIM_NET_59));

   NOT_GATE      GATE_36 (.Input_1(s_LOGISIM_NET_17),
                          .Result(s_LOGISIM_NET_501));

   NOT_GATE      GATE_37 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_772));

   NOT_GATE      GATE_38 (.Input_1(s_LOGISIM_NET_17),
                          .Result(s_LOGISIM_NET_485));

   NOT_GATE      GATE_39 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_750));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_40 (.Input_1(s_LOGISIM_NET_7),
               .Input_2(s_LOGISIM_NET_9),
               .Input_3(s_LOGISIM_NET_8),
               .Input_4(s_LOGISIM_NET_802),
               .Input_5(s_LOGISIM_NET_386),
               .Input_6(s_LOGISIM_NET_3),
               .Input_7(s_LOGISIM_NET_280),
               .Input_8(s_LOGISIM_NET_74),
               .Result(s_LOGISIM_NET_316));

   NOT_GATE      GATE_41 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_620));

   NOT_GATE      GATE_42 (.Input_1(s_LOGISIM_NET_54),
                          .Result(s_LOGISIM_NET_248));

   NOT_GATE      GATE_43 (.Input_1(s_LOGISIM_NET_54),
                          .Result(s_LOGISIM_NET_803));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_44 (.Input_1(s_LOGISIM_NET_7),
               .Input_2(s_LOGISIM_NET_307),
               .Input_3(s_LOGISIM_NET_8),
               .Input_4(s_LOGISIM_NET_759),
               .Input_5(s_LOGISIM_NET_306),
               .Input_6(s_LOGISIM_NET_401),
               .Input_7(s_LOGISIM_NET_631),
               .Input_8(s_LOGISIM_NET_263),
               .Result(s_LOGISIM_NET_703));

   NOT_GATE      GATE_45 (.Input_1(s_LOGISIM_NET_54),
                          .Result(s_LOGISIM_NET_41));

   NOT_GATE      GATE_46 (.Input_1(s_LOGISIM_NET_10),
                          .Result(s_LOGISIM_NET_33));

   NOT_GATE      GATE_47 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_67));

   NOT_GATE      GATE_48 (.Input_1(s_LOGISIM_NET_10),
                          .Result(s_LOGISIM_NET_603));

   NOT_GATE      GATE_49 (.Input_1(s_LOGISIM_NET_3),
                          .Result(s_LOGISIM_NET_477));

   NOT_GATE      GATE_50 (.Input_1(s_LOGISIM_NET_17),
                          .Result(s_LOGISIM_NET_228));

   NOT_GATE      GATE_51 (.Input_1(s_LOGISIM_NET_21),
                          .Result(s_LOGISIM_NET_16));

   NOT_GATE      GATE_52 (.Input_1(s_LOGISIM_NET_9),
                          .Result(s_LOGISIM_NET_755));

   NOT_GATE      GATE_53 (.Input_1(s_LOGISIM_NET_10),
                          .Result(s_LOGISIM_NET_337));

   NOT_GATE      GATE_54 (.Input_1(s_LOGISIM_NET_17),
                          .Result(s_LOGISIM_NET_530));

   NOT_GATE      GATE_55 (.Input_1(s_LOGISIM_NET_54),
                          .Result(s_LOGISIM_NET_494));

   NOT_GATE      GATE_56 (.Input_1(s_LOGISIM_NET_21),
                          .Result(s_LOGISIM_NET_112));

   OR_GATE #(.BubblesMask(0))
      GATE_57 (.Input_1(s_LOGISIM_NET_273),
               .Input_2(s_LOGISIM_NET_794),
               .Result(s_LOGISIM_NET_670));

   NOT_GATE      GATE_58 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_741));

   NOT_GATE      GATE_59 (.Input_1(s_LOGISIM_NET_17),
                          .Result(s_LOGISIM_NET_524));

   NOT_GATE      GATE_60 (.Input_1(s_LOGISIM_NET_54),
                          .Result(s_LOGISIM_NET_216));

   NOT_GATE      GATE_61 (.Input_1(s_LOGISIM_NET_17),
                          .Result(s_LOGISIM_NET_671));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_62 (.Input_1(s_LOGISIM_NET_545),
               .Input_10(s_LOGISIM_NET_228),
               .Input_2(s_LOGISIM_NET_495),
               .Input_3(s_LOGISIM_NET_393),
               .Input_4(s_LOGISIM_NET_253),
               .Input_5(s_LOGISIM_NET_793),
               .Input_6(s_LOGISIM_NET_216),
               .Input_7(s_LOGISIM_NET_21),
               .Input_8(s_LOGISIM_NET_3),
               .Input_9(s_LOGISIM_NET_218),
               .Result(s_LOGISIM_NET_584));

   NOT_GATE      GATE_63 (.Input_1(s_LOGISIM_NET_17),
                          .Result(s_LOGISIM_NET_390));

   NOT_GATE      GATE_64 (.Input_1(s_LOGISIM_NET_20),
                          .Result(s_LOGISIM_NET_203));

   NOT_GATE      GATE_65 (.Input_1(s_LOGISIM_NET_17),
                          .Result(s_LOGISIM_NET_159));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_66 (.Input_1(s_LOGISIM_NET_7),
               .Input_2(s_LOGISIM_NET_428),
               .Input_3(s_LOGISIM_NET_304),
               .Input_4(s_LOGISIM_NET_54),
               .Input_5(s_LOGISIM_NET_21),
               .Input_6(s_LOGISIM_NET_536),
               .Input_7(s_LOGISIM_NET_48),
               .Input_8(s_LOGISIM_NET_342),
               .Result(s_LOGISIM_NET_220));

   NOT_GATE      GATE_67 (.Input_1(s_LOGISIM_NET_20),
                          .Result(s_LOGISIM_NET_278));

   NOT_GATE      GATE_68 (.Input_1(s_LOGISIM_NET_3),
                          .Result(s_LOGISIM_NET_58));

   NOT_GATE      GATE_69 (.Input_1(s_LOGISIM_NET_10),
                          .Result(s_LOGISIM_NET_445));

   NOT_GATE      GATE_70 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_564));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_71 (.Input_1(s_LOGISIM_NET_689),
               .Input_10(s_LOGISIM_NET_490),
               .Input_2(s_LOGISIM_NET_658),
               .Input_3(s_LOGISIM_NET_591),
               .Input_4(s_LOGISIM_NET_511),
               .Input_5(s_LOGISIM_NET_227),
               .Input_6(s_LOGISIM_NET_54),
               .Input_7(s_LOGISIM_NET_21),
               .Input_8(s_LOGISIM_NET_3),
               .Input_9(s_LOGISIM_NET_111),
               .Result(s_LOGISIM_NET_804));

   NOT_GATE      GATE_72 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_246));

   NOT_GATE      GATE_73 (.Input_1(s_LOGISIM_NET_21),
                          .Result(s_LOGISIM_NET_375));

   OR_GATE #(.BubblesMask(0))
      GATE_74 (.Input_1(s_LOGISIM_NET_267),
               .Input_2(s_LOGISIM_NET_683),
               .Result(s_LOGISIM_NET_324));

   NOT_GATE      GATE_75 (.Input_1(s_LOGISIM_NET_54),
                          .Result(s_LOGISIM_NET_417));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_76 (.Input_1(s_LOGISIM_NET_367),
               .Input_10(s_LOGISIM_NET_665),
               .Input_2(s_LOGISIM_NET_140),
               .Input_3(s_LOGISIM_NET_100),
               .Input_4(s_LOGISIM_NET_9),
               .Input_5(s_LOGISIM_NET_8),
               .Input_6(s_LOGISIM_NET_579),
               .Input_7(s_LOGISIM_NET_21),
               .Input_8(s_LOGISIM_NET_3),
               .Input_9(s_LOGISIM_NET_446),
               .Result(s_LOGISIM_NET_756));

   NOT_GATE      GATE_77 (.Input_1(s_LOGISIM_NET_10),
                          .Result(s_LOGISIM_NET_590));

   NOT_GATE      GATE_78 (.Input_1(s_LOGISIM_NET_8),
                          .Result(s_LOGISIM_NET_644));

   NOT_GATE      GATE_79 (.Input_1(s_LOGISIM_NET_10),
                          .Result(s_LOGISIM_NET_32));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_80 (.Input_1(s_LOGISIM_NET_624),
               .Input_10(s_LOGISIM_NET_330),
               .Input_2(s_LOGISIM_NET_586),
               .Input_3(s_LOGISIM_NET_499),
               .Input_4(s_LOGISIM_NET_399),
               .Input_5(s_LOGISIM_NET_8),
               .Input_6(s_LOGISIM_NET_54),
               .Input_7(s_LOGISIM_NET_587),
               .Input_8(s_LOGISIM_NET_3),
               .Input_9(s_LOGISIM_NET_57),
               .Result(s_LOGISIM_NET_787));

   NOT_GATE      GATE_81 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_654));

   NOT_GATE      GATE_82 (.Input_1(s_LOGISIM_NET_3),
                          .Result(s_LOGISIM_NET_185));

   NOT_GATE      GATE_83 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_626));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_84 (.Input_1(s_LOGISIM_NET_592),
               .Input_2(s_LOGISIM_NET_510),
               .Input_3(s_LOGISIM_NET_54),
               .Input_4(s_LOGISIM_NET_150),
               .Input_5(s_LOGISIM_NET_3),
               .Input_6(s_LOGISIM_NET_245),
               .Input_7(s_LOGISIM_NET_444),
               .Result(s_LOGISIM_NET_733));

   NOT_GATE      GATE_85 (.Input_1(s_LOGISIM_NET_9),
                          .Result(s_LOGISIM_NET_160));

   NOT_GATE      GATE_86 (.Input_1(s_LOGISIM_NET_17),
                          .Result(s_LOGISIM_NET_351));

   NOT_GATE      GATE_87 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_408));

   NOT_GATE      GATE_88 (.Input_1(s_LOGISIM_NET_21),
                          .Result(s_LOGISIM_NET_622));

   NOT_GATE      GATE_89 (.Input_1(s_LOGISIM_NET_54),
                          .Result(s_LOGISIM_NET_329));

   NOT_GATE      GATE_90 (.Input_1(s_LOGISIM_NET_8),
                          .Result(s_LOGISIM_NET_356));

   NOT_GATE      GATE_91 (.Input_1(s_LOGISIM_NET_10),
                          .Result(s_LOGISIM_NET_82));

   NOT_GATE      GATE_92 (.Input_1(s_LOGISIM_NET_8),
                          .Result(s_LOGISIM_NET_193));

   NOT_GATE      GATE_93 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_727));

   NOT_GATE      GATE_94 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_269));

   NOT_GATE      GATE_95 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_555));

   NOT_GATE      GATE_96 (.Input_1(s_LOGISIM_NET_17),
                          .Result(s_LOGISIM_NET_583));

   NOT_GATE      GATE_97 (.Input_1(s_LOGISIM_NET_8),
                          .Result(s_LOGISIM_NET_312));

   NOT_GATE      GATE_98 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_641));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_99 (.Input_1(s_LOGISIM_NET_103),
               .Input_10(s_LOGISIM_NET_559),
               .Input_2(s_LOGISIM_NET_735),
               .Input_3(s_LOGISIM_NET_687),
               .Input_4(s_LOGISIM_NET_9),
               .Input_5(s_LOGISIM_NET_328),
               .Input_6(s_LOGISIM_NET_120),
               .Input_7(s_LOGISIM_NET_21),
               .Input_8(s_LOGISIM_NET_3),
               .Input_9(s_LOGISIM_NET_252),
               .Result(s_LOGISIM_NET_567));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_100 (.Input_1(s_LOGISIM_NET_231),
                .Input_10(s_LOGISIM_NET_761),
                .Input_2(s_LOGISIM_NET_118),
                .Input_3(s_LOGISIM_NET_7),
                .Input_4(s_LOGISIM_NET_25),
                .Input_5(s_LOGISIM_NET_8),
                .Input_6(s_LOGISIM_NET_719),
                .Input_7(s_LOGISIM_NET_333),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_638),
                .Result(s_LOGISIM_NET_55));

   NOT_GATE      GATE_101 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_698));

   NOT_GATE      GATE_102 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_535));

   NOT_GATE      GATE_103 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_438));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_104 (.Input_1(s_LOGISIM_NET_20),
                .Input_10(s_LOGISIM_NET_93),
                .Input_2(s_LOGISIM_NET_425),
                .Input_3(s_LOGISIM_NET_302),
                .Input_4(s_LOGISIM_NET_119),
                .Input_5(s_LOGISIM_NET_785),
                .Input_6(s_LOGISIM_NET_79),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_82),
                .Result(s_LOGISIM_NET_338));

   NOT_GATE      GATE_105 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_152));

   NOT_GATE      GATE_106 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_101));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_107 (.Input_1(s_LOGISIM_NET_652),
                .Input_10(s_LOGISIM_NET_385),
                .Input_2(s_LOGISIM_NET_616),
                .Input_3(s_LOGISIM_NET_539),
                .Input_4(s_LOGISIM_NET_432),
                .Input_5(s_LOGISIM_NET_8),
                .Input_6(s_LOGISIM_NET_186),
                .Input_7(s_LOGISIM_NET_16),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_141),
                .Result(s_LOGISIM_NET_389));

   NOT_GATE      GATE_108 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_424));

   NOT_GATE      GATE_109 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_678));

   NOT_GATE      GATE_110 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_261));

   NOT_GATE      GATE_111 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_250));

   NOT_GATE      GATE_112 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_330));

   NOT_GATE      GATE_113 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_690));

   NOT_GATE      GATE_114 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_742));

   NOT_GATE      GATE_115 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_495));

   NOT_GATE      GATE_116 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_368));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_117 (.Input_1(s_LOGISIM_NET_322),
                .Input_2(s_LOGISIM_NET_76),
                .Input_3(s_LOGISIM_NET_54),
                .Input_4(s_LOGISIM_NET_709),
                .Input_5(s_LOGISIM_NET_3),
                .Input_6(s_LOGISIM_NET_179),
                .Input_7(s_LOGISIM_NET_520),
                .Result(s_LOGISIM_NET_472));

   NOT_GATE      GATE_118 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_238));

   NOT_GATE      GATE_119 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_528));

   NOT_GATE      GATE_120 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_215));

   NOT_GATE      GATE_121 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_111));

   NOT_GATE      GATE_122 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_385));

   NOT_GATE      GATE_123 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_720));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_124 (.Input_1(s_LOGISIM_NET_649),
                .Input_2(s_LOGISIM_NET_581),
                .Input_3(s_LOGISIM_NET_486),
                .Input_4(s_LOGISIM_NET_54),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_35),
                .Input_7(s_LOGISIM_NET_336),
                .Input_8(s_LOGISIM_NET_17),
                .Result(s_LOGISIM_NET_264));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_125 (.Input_1(s_LOGISIM_NET_751),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_597),
                .Input_4(s_LOGISIM_NET_331),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_340),
                .Input_7(s_LOGISIM_NET_33),
                .Input_8(s_LOGISIM_NET_315),
                .Result(s_LOGISIM_NET_273));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_126 (.Input_1(s_LOGISIM_NET_380),
                .Input_10(s_LOGISIM_NET_671),
                .Input_2(s_LOGISIM_NET_161),
                .Input_3(s_LOGISIM_NET_744),
                .Input_4(s_LOGISIM_NET_125),
                .Input_5(s_LOGISIM_NET_8),
                .Input_6(s_LOGISIM_NET_54),
                .Input_7(s_LOGISIM_NET_475),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_455),
                .Result(s_LOGISIM_NET_397));

   NOT_GATE      GATE_127 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_486));

   NOT_GATE      GATE_128 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_553));

   NOT_GATE      GATE_129 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_106));

   NOT_GATE      GATE_130 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_376));

   NOT_GATE      GATE_131 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_487));

   NOT_GATE      GATE_132 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_661));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_133 (.Input_1(s_LOGISIM_NET_457),
                .Input_2(s_LOGISIM_NET_348),
                .Input_3(s_LOGISIM_NET_54),
                .Input_4(s_LOGISIM_NET_798),
                .Input_5(s_LOGISIM_NET_3),
                .Input_6(s_LOGISIM_NET_590),
                .Input_7(s_LOGISIM_NET_266),
                .Result(s_LOGISIM_NET_30));

   NOT_GATE      GATE_134 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_392));

   NOT_GATE      GATE_135 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_120));

   NOT_GATE      GATE_136 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_181));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_137 (.Input_1(s_LOGISIM_NET_270),
                .Input_10(s_LOGISIM_NET_617),
                .Input_2(s_LOGISIM_NET_758),
                .Input_3(s_LOGISIM_NET_7),
                .Input_4(s_LOGISIM_NET_627),
                .Input_5(s_LOGISIM_NET_426),
                .Input_6(s_LOGISIM_NET_282),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_363),
                .Result(s_LOGISIM_NET_593));

   NOT_GATE      GATE_138 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_601));

   NOT_GATE      GATE_139 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_357));

   NOT_GATE      GATE_140 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_650));

   NOT_GATE      GATE_141 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_645));

   NOT_GATE      GATE_142 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_52));

   NOT_GATE      GATE_143 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_225));

   NOT_GATE      GATE_144 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_194));

   NOT_GATE      GATE_145 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_411));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_146 (.Input_1(s_LOGISIM_NET_102),
                .Input_2(s_LOGISIM_NET_384),
                .Input_3(s_LOGISIM_NET_54),
                .Input_4(s_LOGISIM_NET_634),
                .Input_5(s_LOGISIM_NET_3),
                .Input_6(s_LOGISIM_NET_162),
                .Input_7(s_LOGISIM_NET_395),
                .Result(s_LOGISIM_NET_474));

   NOT_GATE      GATE_147 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_197));

   NOT_GATE      GATE_148 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_12));

   NOT_GATE      GATE_149 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_432));

   NOT_GATE      GATE_150 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_299));

   NOT_GATE      GATE_151 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_679));

   NOT_GATE      GATE_152 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_770));

   NOT_GATE      GATE_153 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_580));

   NOT_GATE      GATE_154 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_490));

   NOT_GATE      GATE_155 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_183));

   NOT_GATE      GATE_156 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_542));

   NOT_GATE      GATE_157 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_234));

   NOT_GATE      GATE_158 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_282));

   NOT_GATE      GATE_159 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_214));

   NOT_GATE      GATE_160 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_447));

   NOT_GATE      GATE_161 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_180));

   AND_GATE_5_INPUTS #(.BubblesMask(0))
      GATE_162 (.Input_1(s_LOGISIM_NET_544),
                .Input_2(s_LOGISIM_NET_21),
                .Input_3(s_LOGISIM_NET_3),
                .Input_4(s_LOGISIM_NET_487),
                .Input_5(s_LOGISIM_NET_17),
                .Result(s_LOGISIM_NET_561));

   NOT_GATE      GATE_163 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_283));

   NOT_GATE      GATE_164 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_259));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_165 (.Input_1(s_LOGISIM_NET_59),
                .Input_2(s_LOGISIM_NET_260),
                .Input_3(s_LOGISIM_NET_54),
                .Input_4(s_LOGISIM_NET_748),
                .Input_5(s_LOGISIM_NET_3),
                .Input_6(s_LOGISIM_NET_317),
                .Input_7(s_LOGISIM_NET_594),
                .Result(s_LOGISIM_NET_325));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_166 (.Input_1(s_LOGISIM_NET_7),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_213),
                .Input_4(s_LOGISIM_NET_54),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_3),
                .Input_7(s_LOGISIM_NET_130),
                .Input_8(s_LOGISIM_NET_498),
                .Result(s_LOGISIM_NET_175));

   NOT_GATE      GATE_167 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_123));

   NOT_GATE      GATE_168 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_702));

   NOT_GATE      GATE_169 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_147));

   NOT_GATE      GATE_170 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_668));

   NOT_GATE      GATE_171 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_395));

   NOT_GATE      GATE_172 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_480));

   NOT_GATE      GATE_173 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_414));

   NOT_GATE      GATE_174 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_230));

   NOT_GATE      GATE_175 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_722));

   NOT_GATE      GATE_176 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_716));

   NOT_GATE      GATE_177 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_550));

   NOT_GATE      GATE_178 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_363));

   NOT_GATE      GATE_179 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_457));

   NOT_GATE      GATE_180 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_237));

   NOT_GATE      GATE_181 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_585));

   NOT_GATE      GATE_182 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_263));

   NOT_GATE      GATE_183 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_307));

   NOT_GATE      GATE_184 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_87));

   NOT_GATE      GATE_185 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_768));

   NOT_GATE      GATE_186 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_461));

   NOT_GATE      GATE_187 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_353));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_188 (.Input_1(s_LOGISIM_NET_277),
                .Input_2(s_LOGISIM_NET_67),
                .Input_3(s_LOGISIM_NET_54),
                .Input_4(s_LOGISIM_NET_770),
                .Input_5(s_LOGISIM_NET_3),
                .Input_6(s_LOGISIM_NET_440),
                .Input_7(s_LOGISIM_NET_666),
                .Result(s_LOGISIM_NET_339));

   NOT_GATE      GATE_189 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_471));

   NOT_GATE      GATE_190 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_687));

   NOT_GATE      GATE_191 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_536));

   NOT_GATE      GATE_192 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_103));

   NOT_GATE      GATE_193 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_409));

   NOT_GATE      GATE_194 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_245));

   NOT_GATE      GATE_195 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_667));

   NOT_GATE      GATE_196 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_384));

   NOT_GATE      GATE_197 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_360));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_198 (.Input_1(s_LOGISIM_NET_258),
                .Input_2(s_LOGISIM_NET_51),
                .Input_3(s_LOGISIM_NET_54),
                .Input_4(s_LOGISIM_NET_768),
                .Input_5(s_LOGISIM_NET_3),
                .Input_6(s_LOGISIM_NET_435),
                .Input_7(s_LOGISIM_NET_657),
                .Result(s_LOGISIM_NET_436));

   NOT_GATE      GATE_199 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_266));

   NOT_GATE      GATE_200 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_310));

   NOT_GATE      GATE_201 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_718));

   OR_GATE_14_INPUTS #(.BubblesMask(0))
      GATE_202 (.Input_1(s_LOGISIM_NET_275),
                .Input_10(s_LOGISIM_NET_97),
                .Input_11(s_LOGISIM_NET_344),
                .Input_12(s_LOGISIM_NET_703),
                .Input_13(s_LOGISIM_NET_762),
                .Input_14(s_LOGISIM_NET_122),
                .Input_2(s_LOGISIM_NET_133),
                .Input_3(s_LOGISIM_NET_422),
                .Input_4(s_LOGISIM_NET_184),
                .Input_5(s_LOGISIM_NET_725),
                .Input_6(s_LOGISIM_NET_517),
                .Input_7(s_LOGISIM_NET_55),
                .Input_8(s_LOGISIM_NET_646),
                .Input_9(s_LOGISIM_NET_598),
                .Result(s_LOGISIM_NET_226));

   NOT_GATE      GATE_203 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_416));

   NOT_GATE      GATE_204 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_719));

   NOT_GATE      GATE_205 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_170));

   NOT_GATE      GATE_206 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_643));

   NOT_GATE      GATE_207 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_4));

   NOT_GATE      GATE_208 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_623));

   NOT_GATE      GATE_209 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_171));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_210 (.Input_1(s_LOGISIM_NET_525),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_155),
                .Input_4(s_LOGISIM_NET_776),
                .Input_5(s_LOGISIM_NET_112),
                .Input_6(s_LOGISIM_NET_489),
                .Input_7(s_LOGISIM_NET_116),
                .Input_8(s_LOGISIM_NET_17),
                .Result(s_LOGISIM_NET_305));

   NOT_GATE      GATE_211 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_254));

   NOT_GATE      GATE_212 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_642));

   NOT_GATE      GATE_213 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_311));

   NOT_GATE      GATE_214 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_640));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_215 (.Input_1(s_LOGISIM_NET_565),
                .Input_10(s_LOGISIM_NET_107),
                .Input_2(s_LOGISIM_NET_519),
                .Input_3(s_LOGISIM_NET_7),
                .Input_4(s_LOGISIM_NET_137),
                .Input_5(s_LOGISIM_NET_786),
                .Input_6(s_LOGISIM_NET_94),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_95),
                .Result(s_LOGISIM_NET_223));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_216 (.Input_1(s_LOGISIM_NET_482),
                .Input_10(s_LOGISIM_NET_722),
                .Input_2(s_LOGISIM_NET_69),
                .Input_3(s_LOGISIM_NET_71),
                .Input_4(s_LOGISIM_NET_9),
                .Input_5(s_LOGISIM_NET_595),
                .Input_6(s_LOGISIM_NET_494),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_556),
                .Result(s_LOGISIM_NET_85));

   NOT_GATE      GATE_217 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_131));

   NOT_GATE      GATE_218 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_516));

   NOT_GATE      GATE_219 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_427));

   NOT_GATE      GATE_220 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_707));

   NOT_GATE      GATE_221 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_298));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_222 (.Input_1(s_LOGISIM_NET_278),
                .Input_10(s_LOGISIM_NET_614),
                .Input_2(s_LOGISIM_NET_753),
                .Input_3(s_LOGISIM_NET_710),
                .Input_4(s_LOGISIM_NET_650),
                .Input_5(s_LOGISIM_NET_8),
                .Input_6(s_LOGISIM_NET_54),
                .Input_7(s_LOGISIM_NET_396),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_365),
                .Result(s_LOGISIM_NET_145));

   NOT_GATE      GATE_223 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_382));

   NOT_GATE      GATE_224 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_701));

   NOT_GATE      GATE_225 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_597));

   NOT_GATE      GATE_226 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_659));

   NOT_GATE      GATE_227 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_29));

   NOT_GATE      GATE_228 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_281));

   NOT_GATE      GATE_229 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_86));

   NOT_GATE      GATE_230 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_270));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_231 (.Input_1(s_LOGISIM_NET_656),
                .Input_2(s_LOGISIM_NET_589),
                .Input_3(s_LOGISIM_NET_54),
                .Input_4(s_LOGISIM_NET_318),
                .Input_5(s_LOGISIM_NET_3),
                .Input_6(s_LOGISIM_NET_383),
                .Input_7(s_LOGISIM_NET_549),
                .Result(s_LOGISIM_NET_113));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_232 (.Input_1(s_LOGISIM_NET_203),
                .Input_10(s_LOGISIM_NET_774),
                .Input_2(s_LOGISIM_NET_92),
                .Input_3(s_LOGISIM_NET_392),
                .Input_4(s_LOGISIM_NET_171),
                .Input_5(s_LOGISIM_NET_8),
                .Input_6(s_LOGISIM_NET_746),
                .Input_7(s_LOGISIM_NET_98),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_685),
                .Result(s_LOGISIM_NET_517));

   NOT_GATE      GATE_233 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_575));

   NOT_GATE      GATE_234 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_28));

   NOT_GATE      GATE_235 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_591));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_236 (.Input_1(s_LOGISIM_NET_75),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_34),
                .Input_4(s_LOGISIM_NET_468),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_473),
                .Input_7(s_LOGISIM_NET_49),
                .Input_8(s_LOGISIM_NET_460),
                .Result(s_LOGISIM_NET_97));

   NOT_GATE      GATE_237 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_526));

   NOT_GATE      GATE_238 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_469));

   NOT_GATE      GATE_239 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_566));

   NOT_GATE      GATE_240 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_574));

   NOT_GATE      GATE_241 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_430));

   NOT_GATE      GATE_242 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_213));

   NOT_GATE      GATE_243 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_361));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_244 (.Input_1(s_LOGISIM_NET_521),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_138),
                .Input_4(s_LOGISIM_NET_775),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_477),
                .Input_7(s_LOGISIM_NET_680),
                .Input_8(s_LOGISIM_NET_262),
                .Result(s_LOGISIM_NET_267));

   NOT_GATE      GATE_245 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_682));

   NOT_GATE      GATE_246 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_313));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_247 (.Input_1(s_LOGISIM_NET_469),
                .Input_10(s_LOGISIM_NET_64),
                .Input_2(s_LOGISIM_NET_414),
                .Input_3(s_LOGISIM_NET_7),
                .Input_4(s_LOGISIM_NET_9),
                .Input_5(s_LOGISIM_NET_747),
                .Input_6(s_LOGISIM_NET_215),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_724),
                .Result(s_LOGISIM_NET_65));

   NOT_GATE      GATE_248 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_466));

   NOT_GATE      GATE_249 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_506));

   NOT_GATE      GATE_250 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_521));

   NOT_GATE      GATE_251 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_587));

   NOT_GATE      GATE_252 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_61));

   NOT_GATE      GATE_253 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_401));

   NOT_GATE      GATE_254 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_127));

   NOT_GATE      GATE_255 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_773));

   NOT_GATE      GATE_256 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_129));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_257 (.Input_1(s_LOGISIM_NET_7),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_8),
                .Input_4(s_LOGISIM_NET_692),
                .Input_5(s_LOGISIM_NET_647),
                .Input_6(s_LOGISIM_NET_3),
                .Input_7(s_LOGISIM_NET_492),
                .Input_8(s_LOGISIM_NET_688),
                .Result(s_LOGISIM_NET_133));

   NOT_GATE      GATE_258 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_404));

   NOT_GATE      GATE_259 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_450));

   NOT_GATE      GATE_260 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_380));

   NOT_GATE      GATE_261 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_511));

   NOT_GATE      GATE_262 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_637));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_263 (.Input_1(s_LOGISIM_NET_607),
                .Input_10(s_LOGISIM_NET_298),
                .Input_2(s_LOGISIM_NET_571),
                .Input_3(s_LOGISIM_NET_471),
                .Input_4(s_LOGISIM_NET_361),
                .Input_5(s_LOGISIM_NET_8),
                .Input_6(s_LOGISIM_NET_54),
                .Input_7(s_LOGISIM_NET_574),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_285),
                .Result(s_LOGISIM_NET_165));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_264 (.Input_1(s_LOGISIM_NET_562),
                .Input_10(s_LOGISIM_NET_754),
                .Input_2(s_LOGISIM_NET_66),
                .Input_3(s_LOGISIM_NET_237),
                .Input_4(s_LOGISIM_NET_357),
                .Input_5(s_LOGISIM_NET_648),
                .Input_6(s_LOGISIM_NET_54),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_611),
                .Result(s_LOGISIM_NET_636));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_265 (.Input_1(s_LOGISIM_NET_661),
                .Input_10(s_LOGISIM_NET_295),
                .Input_2(s_LOGISIM_NET_626),
                .Input_3(s_LOGISIM_NET_7),
                .Input_4(s_LOGISIM_NET_360),
                .Input_5(s_LOGISIM_NET_8),
                .Input_6(s_LOGISIM_NET_41),
                .Input_7(s_LOGISIM_NET_578),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_343),
                .Result(s_LOGISIM_NET_247));

   NOT_GATE      GATE_266 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_509));

   NOT_GATE      GATE_267 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_612));

   NOT_GATE      GATE_268 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_751));

   NOT_GATE      GATE_269 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_399));

   NOT_GATE      GATE_270 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_99));

   NOT_GATE      GATE_271 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_433));

   NOT_GATE      GATE_272 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_98));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_273 (.Input_1(s_LOGISIM_NET_7),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_8),
                .Input_4(s_LOGISIM_NET_329),
                .Input_5(s_LOGISIM_NET_210),
                .Input_6(s_LOGISIM_NET_3),
                .Input_7(s_LOGISIM_NET_32),
                .Input_8(s_LOGISIM_NET_314),
                .Result(s_LOGISIM_NET_373));

   NOT_GATE      GATE_274 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_673));

   NOT_GATE      GATE_275 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_410));

   NOT_GATE      GATE_276 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_27));

   NOT_GATE      GATE_277 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_257));

   NOT_GATE      GATE_278 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_431));

   NOT_GATE      GATE_279 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_211));

   NOT_GATE      GATE_280 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_251));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_281 (.Input_1(s_LOGISIM_NET_7),
                .Input_2(s_LOGISIM_NET_535),
                .Input_3(s_LOGISIM_NET_8),
                .Input_4(s_LOGISIM_NET_54),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_560),
                .Input_7(s_LOGISIM_NET_99),
                .Input_8(s_LOGISIM_NET_374),
                .Result(s_LOGISIM_NET_730));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_282 (.Input_1(s_LOGISIM_NET_645),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_405),
                .Input_4(s_LOGISIM_NET_803),
                .Input_5(s_LOGISIM_NET_387),
                .Input_6(s_LOGISIM_NET_124),
                .Input_7(s_LOGISIM_NET_388),
                .Input_8(s_LOGISIM_NET_17),
                .Result(s_LOGISIM_NET_415));

   NOT_GATE      GATE_283 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_318));

   NOT_GATE      GATE_284 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_218));

   NOT_GATE      GATE_285 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_781));

   NOT_GATE      GATE_286 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_610));

   NOT_GATE      GATE_287 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_2));

   NOT_GATE      GATE_288 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_142));

   AND_GATE_5_INPUTS #(.BubblesMask(0))
      GATE_289 (.Input_1(s_LOGISIM_NET_54),
                .Input_2(s_LOGISIM_NET_21),
                .Input_3(s_LOGISIM_NET_516),
                .Input_4(s_LOGISIM_NET_10),
                .Input_5(s_LOGISIM_NET_17),
                .Result(s_LOGISIM_NET_769));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_290 (.Input_1(s_LOGISIM_NET_7),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_268),
                .Input_4(s_LOGISIM_NET_789),
                .Input_5(s_LOGISIM_NET_235),
                .Input_6(s_LOGISIM_NET_3),
                .Input_7(s_LOGISIM_NET_73),
                .Input_8(s_LOGISIM_NET_353),
                .Result(s_LOGISIM_NET_547));

   NOT_GATE      GATE_291 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_138));

   NOT_GATE      GATE_292 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_202));

   NOT_GATE      GATE_293 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_272));

   NOT_GATE      GATE_294 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_473));

   NOT_GATE      GATE_295 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_405));

   NOT_GATE      GATE_296 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_240));

   NOT_GATE      GATE_297 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_364));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_298 (.Input_1(s_LOGISIM_NET_362),
                .Input_10(s_LOGISIM_NET_27),
                .Input_2(s_LOGISIM_NET_290),
                .Input_3(s_LOGISIM_NET_7),
                .Input_4(s_LOGISIM_NET_286),
                .Input_5(s_LOGISIM_NET_742),
                .Input_6(s_LOGISIM_NET_191),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_716),
                .Result(s_LOGISIM_NET_697));

   NOT_GATE      GATE_299 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_426));

   NOT_GATE      GATE_300 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_546));

   NOT_GATE      GATE_301 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_221));

   NOT_GATE      GATE_302 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_565));

   OR_GATE_17_INPUTS #(.BubblesMask(0))
      GATE_303 (.Input_1(s_LOGISIM_NET_105),
                .Input_10(s_LOGISIM_NET_296),
                .Input_11(s_LOGISIM_NET_593),
                .Input_12(s_LOGISIM_NET_309),
                .Input_13(s_LOGISIM_NET_220),
                .Input_14(s_LOGISIM_NET_421),
                .Input_15(s_LOGISIM_NET_663),
                .Input_16(s_LOGISIM_NET_633),
                .Input_17(s_LOGISIM_NET_113),
                .Input_2(s_LOGISIM_NET_358),
                .Input_3(s_LOGISIM_NET_117),
                .Input_4(s_LOGISIM_NET_660),
                .Input_5(s_LOGISIM_NET_567),
                .Input_6(s_LOGISIM_NET_88),
                .Input_7(s_LOGISIM_NET_37),
                .Input_8(s_LOGISIM_NET_514),
                .Input_9(s_LOGISIM_NET_178),
                .Result(s_LOGISIM_NET_795));

   NOT_GATE      GATE_304 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_448));

   NOT_GATE      GATE_305 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_374));

   NOT_GATE      GATE_306 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_104));

   NOT_GATE      GATE_307 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_412));

   NOT_GATE      GATE_308 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_570));

   NOT_GATE      GATE_309 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_712));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_310 (.Input_1(s_LOGISIM_NET_570),
                .Input_2(s_LOGISIM_NET_476),
                .Input_3(s_LOGISIM_NET_364),
                .Input_4(s_LOGISIM_NET_800),
                .Input_5(s_LOGISIM_NET_345),
                .Input_6(s_LOGISIM_NET_3),
                .Input_7(s_LOGISIM_NET_222),
                .Input_8(s_LOGISIM_NET_433),
                .Result(s_LOGISIM_NET_275));

   NOT_GATE      GATE_311 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_458));

   NOT_GATE      GATE_312 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_232));

   NOT_GATE      GATE_313 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_478));

   NOT_GATE      GATE_314 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_155));

   NOT_GATE      GATE_315 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_423));

   NOT_GATE      GATE_316 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_572));

   NOT_GATE      GATE_317 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_128));

   NOT_GATE      GATE_318 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_476));

   NOT_GATE      GATE_319 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_749));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_320 (.Input_1(s_LOGISIM_NET_7),
                .Input_2(s_LOGISIM_NET_160),
                .Input_3(s_LOGISIM_NET_356),
                .Input_4(s_LOGISIM_NET_623),
                .Input_5(s_LOGISIM_NET_569),
                .Input_6(s_LOGISIM_NET_3),
                .Input_7(s_LOGISIM_NET_366),
                .Input_8(s_LOGISIM_NET_615),
                .Result(s_LOGISIM_NET_379));

   NOT_GATE      GATE_321 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_695));

   NOT_GATE      GATE_322 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_140));

   NOT_GATE      GATE_323 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_69));

   NOT_GATE      GATE_324 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_757));

   NOT_GATE      GATE_325 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_141));

   NOT_GATE      GATE_326 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_100));

   NOT_GATE      GATE_327 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_456));

   NOT_GATE      GATE_328 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_765));

   NOT_GATE      GATE_329 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_665));

   NOT_GATE      GATE_330 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_792));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_331 (.Input_1(s_LOGISIM_NET_750),
                .Input_2(s_LOGISIM_NET_702),
                .Input_3(s_LOGISIM_NET_640),
                .Input_4(s_LOGISIM_NET_54),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_382),
                .Input_7(s_LOGISIM_NET_104),
                .Input_8(s_LOGISIM_NET_17),
                .Result(s_LOGISIM_NET_40));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_332 (.Input_1(s_LOGISIM_NET_132),
                .Input_10(s_LOGISIM_NET_718),
                .Input_2(s_LOGISIM_NET_4),
                .Input_3(s_LOGISIM_NET_7),
                .Input_4(s_LOGISIM_NET_9),
                .Input_5(s_LOGISIM_NET_8),
                .Input_6(s_LOGISIM_NET_639),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_550),
                .Result(s_LOGISIM_NET_117));

   NOT_GATE      GATE_333 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_25));

   NOT_GATE      GATE_334 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_496));

   NOT_GATE      GATE_335 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_746));

   NOT_GATE      GATE_336 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_462));

   NOT_GATE      GATE_337 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_388));

   NOT_GATE      GATE_338 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_658));

   NOT_GATE      GATE_339 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_761));

   NOT_GATE      GATE_340 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_143));

   NOT_GATE      GATE_341 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_286));

   NOT_GATE      GATE_342 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_497));

   NOT_GATE      GATE_343 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_465));

   NOT_GATE      GATE_344 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_75));

   NOT_GATE      GATE_345 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_95));

   NOT_GATE      GATE_346 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_558));

   OR_GATE_3_INPUTS #(.BubblesMask(0))
      GATE_347 (.Input_1(s_LOGISIM_NET_42),
                .Input_2(s_LOGISIM_NET_784),
                .Input_3(s_LOGISIM_NET_325),
                .Result(s_LOGISIM_NET_766));

   NOT_GATE      GATE_348 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_253));

   NOT_GATE      GATE_349 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_70));

   NOT_GATE      GATE_350 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_607));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_351 (.Input_1(s_LOGISIM_NET_209),
                .Input_2(s_LOGISIM_NET_755),
                .Input_3(s_LOGISIM_NET_183),
                .Input_4(s_LOGISIM_NET_533),
                .Input_5(s_LOGISIM_NET_458),
                .Input_6(s_LOGISIM_NET_3),
                .Input_7(s_LOGISIM_NET_197),
                .Input_8(s_LOGISIM_NET_529),
                .Result(s_LOGISIM_NET_512));

   NOT_GATE      GATE_352 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_508));

   NOT_GATE      GATE_353 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_435));

   NOT_GATE      GATE_354 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_519));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_355 (.Input_1(s_LOGISIM_NET_655),
                .Input_10(s_LOGISIM_NET_127),
                .Input_2(s_LOGISIM_NET_618),
                .Input_3(s_LOGISIM_NET_7),
                .Input_4(s_LOGISIM_NET_9),
                .Input_5(s_LOGISIM_NET_8),
                .Input_6(s_LOGISIM_NET_799),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_23),
                .Result(s_LOGISIM_NET_319));

   NOT_GATE      GATE_356 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_704));

   NOT_GATE      GATE_357 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_710));

   NOT_GATE      GATE_358 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_544));

   NOT_GATE      GATE_359 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_48));

   NOT_GATE      GATE_360 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_758));

   NOT_GATE      GATE_361 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_540));

   NOT_GATE      GATE_362 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_301));

   NOT_GATE      GATE_363 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_31));

   NOT_GATE      GATE_364 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_235));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_365 (.Input_1(s_LOGISIM_NET_189),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_321),
                .Input_4(s_LOGISIM_NET_605),
                .Input_5(s_LOGISIM_NET_553),
                .Input_6(s_LOGISIM_NET_3),
                .Input_7(s_LOGISIM_NET_337),
                .Input_8(s_LOGISIM_NET_600),
                .Result(s_LOGISIM_NET_204));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_366 (.Input_1(s_LOGISIM_NET_621),
                .Input_2(s_LOGISIM_NET_552),
                .Input_3(s_LOGISIM_NET_54),
                .Input_4(s_LOGISIM_NET_234),
                .Input_5(s_LOGISIM_NET_3),
                .Input_6(s_LOGISIM_NET_303),
                .Input_7(s_LOGISIM_NET_491),
                .Result(s_LOGISIM_NET_797));

   NOT_GATE      GATE_367 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_394));

   NOT_GATE      GATE_368 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_672));

   NOT_GATE      GATE_369 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_335));

   NOT_GATE      GATE_370 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_463));

   NOT_GATE      GATE_371 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_336));

   NOT_GATE      GATE_372 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_260));

   NOT_GATE      GATE_373 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_767));

   NOT_GATE      GATE_374 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_90));

   NOT_GATE      GATE_375 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_529));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_376 (.Input_1(s_LOGISIM_NET_7),
                .Input_2(s_LOGISIM_NET_84),
                .Input_3(s_LOGISIM_NET_259),
                .Input_4(s_LOGISIM_NET_54),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_542),
                .Input_7(s_LOGISIM_NET_194),
                .Input_8(s_LOGISIM_NET_530),
                .Result(s_LOGISIM_NET_219));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_377 (.Input_1(s_LOGISIM_NET_157),
                .Input_2(s_LOGISIM_NET_408),
                .Input_3(s_LOGISIM_NET_54),
                .Input_4(s_LOGISIM_NET_651),
                .Input_5(s_LOGISIM_NET_3),
                .Input_6(s_LOGISIM_NET_211),
                .Input_7(s_LOGISIM_NET_416),
                .Result(s_LOGISIM_NET_633));

   NOT_GATE      GATE_378 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_629));

   NOT_GATE      GATE_379 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_647));

   NOT_GATE      GATE_380 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_482));

   NOT_GATE      GATE_381 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_753));

   NOT_GATE      GATE_382 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_177));

   NOT_GATE      GATE_383 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_149));

   NOT_GATE      GATE_384 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_634));

   NOT_GATE      GATE_385 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_543));

   NOT_GATE      GATE_386 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_664));

   NOT_GATE      GATE_387 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_498));

   NOT_GATE      GATE_388 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_56));

   NOT_GATE      GATE_389 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_729));

   NOT_GATE      GATE_390 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_303));

   NOT_GATE      GATE_391 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_96));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_392 (.Input_1(s_LOGISIM_NET_20),
                .Input_10(s_LOGISIM_NET_418),
                .Input_2(s_LOGISIM_NET_610),
                .Input_3(s_LOGISIM_NET_532),
                .Input_4(s_LOGISIM_NET_429),
                .Input_5(s_LOGISIM_NET_77),
                .Input_6(s_LOGISIM_NET_412),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_208),
                .Result(s_LOGISIM_NET_483));

   NOT_GATE      GATE_393 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_407));

   NOT_GATE      GATE_394 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_739));

   NOT_GATE      GATE_395 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_569));

   NOT_GATE      GATE_396 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_802));

   NOT_GATE      GATE_397 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_513));

   NOT_GATE      GATE_398 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_116));

   NOT_GATE      GATE_399 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_599));

   NOT_GATE      GATE_400 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_505));

   NOT_GATE      GATE_401 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_187));

   NOT_GATE      GATE_402 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_23));

   NOT_GATE      GATE_403 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_280));

   NOT_GATE      GATE_404 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_745));

   NOT_GATE      GATE_405 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_460));

   NOT_GATE      GATE_406 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_592));

   NOT_GATE      GATE_407 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_656));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_408 (.Input_1(s_LOGISIM_NET_7),
                .Input_2(s_LOGISIM_NET_448),
                .Input_3(s_LOGISIM_NET_281),
                .Input_4(s_LOGISIM_NET_738),
                .Input_5(s_LOGISIM_NET_170),
                .Input_6(s_LOGISIM_NET_3),
                .Input_7(s_LOGISIM_NET_577),
                .Input_8(s_LOGISIM_NET_731),
                .Result(s_LOGISIM_NET_403));

   NOT_GATE      GATE_409 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_396));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_410 (.Input_1(s_LOGISIM_NET_727),
                .Input_2(s_LOGISIM_NET_674),
                .Input_3(s_LOGISIM_NET_8),
                .Input_4(s_LOGISIM_NET_54),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_185),
                .Input_7(s_LOGISIM_NET_413),
                .Input_8(s_LOGISIM_NET_144),
                .Result(s_LOGISIM_NET_780));

   NOT_GATE      GATE_411 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_635));

   NOT_GATE      GATE_412 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_413));

   NOT_GATE      GATE_413 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_22));

   NOT_GATE      GATE_414 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_196));

   NOT_GATE      GATE_415 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_308));

   NOT_GATE      GATE_416 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_285));

   NOT_GATE      GATE_417 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_200));

   NOT_GATE      GATE_418 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_611));

   NOT_GATE      GATE_419 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_455));

   NOT_GATE      GATE_420 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_788));

   NOT_GATE      GATE_421 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_400));

   NOT_GATE      GATE_422 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_229));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_423 (.Input_1(s_LOGISIM_NET_686),
                .Input_10(s_LOGISIM_NET_485),
                .Input_2(s_LOGISIM_NET_654),
                .Input_3(s_LOGISIM_NET_585),
                .Input_4(s_LOGISIM_NET_500),
                .Input_5(s_LOGISIM_NET_214),
                .Input_6(s_LOGISIM_NET_479),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_101),
                .Result(s_LOGISIM_NET_604));

   NOT_GATE      GATE_424 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_198));

   NOT_GATE      GATE_425 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_345));

   NOT_GATE      GATE_426 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_5));

   NOT_GATE      GATE_427 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_532));

   NOT_GATE      GATE_428 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_119));

   NOT_GATE      GATE_429 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_209));

   NOT_GATE      GATE_430 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_666));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_431 (.Input_1(s_LOGISIM_NET_173),
                .Input_2(s_LOGISIM_NET_284),
                .Input_3(s_LOGISIM_NET_8),
                .Input_4(s_LOGISIM_NET_54),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_5),
                .Input_7(s_LOGISIM_NET_434),
                .Input_8(s_LOGISIM_NET_659),
                .Result(s_LOGISIM_NET_296));

   NOT_GATE      GATE_432 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_79));

   NOT_GATE      GATE_433 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_6));

   OR_GATE_23_INPUTS #(.BubblesMask(0))
      GATE_434 (.Input_1(s_LOGISIM_NET_604),
                .Input_10(s_LOGISIM_NET_403),
                .Input_11(s_LOGISIM_NET_204),
                .Input_12(s_LOGISIM_NET_771),
                .Input_13(s_LOGISIM_NET_332),
                .Input_14(s_LOGISIM_NET_38),
                .Input_15(s_LOGISIM_NET_134),
                .Input_16(s_LOGISIM_NET_691),
                .Input_17(s_LOGISIM_NET_40),
                .Input_18(s_LOGISIM_NET_223),
                .Input_19(s_LOGISIM_NET_561),
                .Input_2(s_LOGISIM_NET_483),
                .Input_20(s_LOGISIM_NET_527),
                .Input_21(s_LOGISIM_NET_415),
                .Input_22(s_LOGISIM_NET_30),
                .Input_23(s_LOGISIM_NET_472),
                .Input_3(s_LOGISIM_NET_319),
                .Input_4(s_LOGISIM_NET_65),
                .Input_5(s_LOGISIM_NET_669),
                .Input_6(s_LOGISIM_NET_350),
                .Input_7(s_LOGISIM_NET_726),
                .Input_8(s_LOGISIM_NET_373),
                .Input_9(s_LOGISIM_NET_547),
                .Result(s_LOGISIM_NET_68));

   NOT_GATE      GATE_435 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_468));

   NOT_GATE      GATE_436 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_205));

   NOT_GATE      GATE_437 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_451));

   NOT_GATE      GATE_438 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_78));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_439 (.Input_1(s_LOGISIM_NET_564),
                .Input_2(s_LOGISIM_NET_464),
                .Input_3(s_LOGISIM_NET_352),
                .Input_4(s_LOGISIM_NET_54),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_566),
                .Input_7(s_LOGISIM_NET_114),
                .Input_8(s_LOGISIM_NET_17),
                .Result(s_LOGISIM_NET_734));

   NOT_GATE      GATE_440 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_35));

   NOT_GATE      GATE_441 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_648));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_442 (.Input_1(s_LOGISIM_NET_763),
                .Input_2(s_LOGISIM_NET_739),
                .Input_3(s_LOGISIM_NET_8),
                .Input_4(s_LOGISIM_NET_54),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_369),
                .Input_7(s_LOGISIM_NET_90),
                .Input_8(s_LOGISIM_NET_351),
                .Result(s_LOGISIM_NET_60));

   NOT_GATE      GATE_443 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_51));

   NOT_GATE      GATE_444 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_632));

   NOT_GATE      GATE_445 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_638));

   NOT_GATE      GATE_446 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_676));

   NOT_GATE      GATE_447 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_369));

   NOT_GATE      GATE_448 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_442));

   NOT_GATE      GATE_449 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_492));

   NOT_GATE      GATE_450 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_443));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_451 (.Input_1(s_LOGISIM_NET_241),
                .Input_10(s_LOGISIM_NET_606),
                .Input_2(s_LOGISIM_NET_772),
                .Input_3(s_LOGISIM_NET_7),
                .Input_4(s_LOGISIM_NET_9),
                .Input_5(s_LOGISIM_NET_411),
                .Input_6(s_LOGISIM_NET_254),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_346),
                .Result(s_LOGISIM_NET_660));

   NOT_GATE      GATE_452 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_239));

   NOT_GATE      GATE_453 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_242));

   NOT_GATE      GATE_454 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_391));

   NOT_GATE      GATE_455 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_39));

   NOT_GATE      GATE_456 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_624));

   AND_GATE_5_INPUTS #(.BubblesMask(0))
      GATE_457 (.Input_1(s_LOGISIM_NET_54),
                .Input_2(s_LOGISIM_NET_21),
                .Input_3(s_LOGISIM_NET_81),
                .Input_4(s_LOGISIM_NET_10),
                .Input_5(s_LOGISIM_NET_17),
                .Result(s_LOGISIM_NET_691));

   NOT_GATE      GATE_458 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_737));

   NOT_GATE      GATE_459 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_752));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_460 (.Input_1(s_LOGISIM_NET_506),
                .Input_10(s_LOGISIM_NET_62),
                .Input_2(s_LOGISIM_NET_452),
                .Input_3(s_LOGISIM_NET_334),
                .Input_4(s_LOGISIM_NET_168),
                .Input_5(s_LOGISIM_NET_8),
                .Input_6(s_LOGISIM_NET_54),
                .Input_7(s_LOGISIM_NET_454),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_43),
                .Result(s_LOGISIM_NET_481));

   NOT_GATE      GATE_461 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_609));

   NOT_GATE      GATE_462 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_110));

   NOT_GATE      GATE_463 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_362));

   NOT_GATE      GATE_464 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_694));

   NOT_GATE      GATE_465 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_428));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_466 (.Input_1(s_LOGISIM_NET_187),
                .Input_10(s_LOGISIM_NET_757),
                .Input_2(s_LOGISIM_NET_72),
                .Input_3(s_LOGISIM_NET_269),
                .Input_4(s_LOGISIM_NET_9),
                .Input_5(s_LOGISIM_NET_8),
                .Input_6(s_LOGISIM_NET_706),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_625),
                .Result(s_LOGISIM_NET_350));

   NOT_GATE      GATE_467 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_531));

   NOT_GATE      GATE_468 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_174));

   NOT_GATE      GATE_469 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_759));

   NOT_GATE      GATE_470 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_439));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_471 (.Input_1(s_LOGISIM_NET_181),
                .Input_2(s_LOGISIM_NET_46),
                .Input_3(s_LOGISIM_NET_225),
                .Input_4(s_LOGISIM_NET_54),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_526),
                .Input_7(s_LOGISIM_NET_154),
                .Input_8(s_LOGISIM_NET_515),
                .Result(s_LOGISIM_NET_192));

   NOT_GATE      GATE_472 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_367));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_473 (.Input_1(s_LOGISIM_NET_7),
                .Input_2(s_LOGISIM_NET_677),
                .Input_3(s_LOGISIM_NET_8),
                .Input_4(s_LOGISIM_NET_248),
                .Input_5(s_LOGISIM_NET_89),
                .Input_6(s_LOGISIM_NET_370),
                .Input_7(s_LOGISIM_NET_538),
                .Input_8(s_LOGISIM_NET_236),
                .Result(s_LOGISIM_NET_527));

   NOT_GATE      GATE_474 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_208));

   NOT_GATE      GATE_475 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_651));

   NOT_GATE      GATE_476 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_446));

   NOT_GATE      GATE_477 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_699));

   NOT_GATE      GATE_478 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_371));

   NOT_GATE      GATE_479 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_57));

   NOT_GATE      GATE_480 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_589));

   NOT_GATE      GATE_481 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_91));

   NOT_GATE      GATE_482 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_13));

   NOT_GATE      GATE_483 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_614));

   NOT_GATE      GATE_484 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_747));

   NOT_GATE      GATE_485 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_608));

   NOT_GATE      GATE_486 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_26));

   NOT_GATE      GATE_487 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_500));

   NOT_GATE      GATE_488 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_53));

   NOT_GATE      GATE_489 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_210));

   NOT_GATE      GATE_490 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_233));

   NOT_GATE      GATE_491 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_686));

   NOT_GATE      GATE_492 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_243));

   NOT_GATE      GATE_493 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_434));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_494 (.Input_1(s_LOGISIM_NET_765),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_643),
                .Input_4(s_LOGISIM_NET_419),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_424),
                .Input_7(s_LOGISIM_NET_202),
                .Input_8(s_LOGISIM_NET_17),
                .Result(s_LOGISIM_NET_372));

   NOT_GATE      GATE_495 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_19));

   NOT_GATE      GATE_496 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_300));

   NOT_GATE      GATE_497 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_782));

   NOT_GATE      GATE_498 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_340));

   NOT_GATE      GATE_499 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_63));

   NOT_GATE      GATE_500 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_464));

   NOT_GATE      GATE_501 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_49));

   NOT_GATE      GATE_502 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_776));

   NOT_GATE      GATE_503 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_92));

   NOT_GATE      GATE_504 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_662));

   NOT_GATE      GATE_505 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_523));

   NOT_GATE      GATE_506 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_588));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_507 (.Input_1(s_LOGISIM_NET_554),
                .Input_2(s_LOGISIM_NET_441),
                .Input_3(s_LOGISIM_NET_54),
                .Input_4(s_LOGISIM_NET_26),
                .Input_5(s_LOGISIM_NET_3),
                .Input_6(s_LOGISIM_NET_126),
                .Input_7(s_LOGISIM_NET_390),
                .Result(s_LOGISIM_NET_784));

   NOT_GATE      GATE_508 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_304));

   NOT_GATE      GATE_509 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_153));

   NOT_GATE      GATE_510 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_552));

   NOT_GATE      GATE_511 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_743));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_512 (.Input_1(s_LOGISIM_NET_299),
                .Input_10(s_LOGISIM_NET_777),
                .Input_2(s_LOGISIM_NET_212),
                .Input_3(s_LOGISIM_NET_406),
                .Input_4(s_LOGISIM_NET_9),
                .Input_5(s_LOGISIM_NET_720),
                .Input_6(s_LOGISIM_NET_78),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_690),
                .Result(s_LOGISIM_NET_669));

   NOT_GATE      GATE_513 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_571));

   NOT_GATE      GATE_514 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_346));

   NOT_GATE      GATE_515 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_347));

   NOT_GATE      GATE_516 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_45));

   NOT_GATE      GATE_517 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_322));

   NOT_GATE      GATE_518 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_596));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_519 (.Input_1(s_LOGISIM_NET_7),
                .Input_2(s_LOGISIM_NET_582),
                .Input_3(s_LOGISIM_NET_488),
                .Input_4(s_LOGISIM_NET_109),
                .Input_5(s_LOGISIM_NET_470),
                .Input_6(s_LOGISIM_NET_3),
                .Input_7(s_LOGISIM_NET_391),
                .Input_8(s_LOGISIM_NET_91),
                .Result(s_LOGISIM_NET_184));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_520 (.Input_1(s_LOGISIM_NET_7),
                .Input_2(s_LOGISIM_NET_196),
                .Input_3(s_LOGISIM_NET_8),
                .Input_4(s_LOGISIM_NET_54),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_513),
                .Input_7(s_LOGISIM_NET_115),
                .Input_8(s_LOGISIM_NET_496),
                .Result(s_LOGISIM_NET_255));

   NOT_GATE      GATE_521 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_327));

   NOT_GATE      GATE_522 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_341));

   NOT_GATE      GATE_523 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_763));

   NOT_GATE      GATE_524 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_774));

   NOT_GATE      GATE_525 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_489));

   NOT_GATE      GATE_526 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_47));

   NOT_GATE      GATE_527 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_291));

   NOT_GATE      GATE_528 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_306));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_529 (.Input_1(s_LOGISIM_NET_180),
                .Input_10(s_LOGISIM_NET_583),
                .Input_2(s_LOGISIM_NET_732),
                .Input_3(s_LOGISIM_NET_681),
                .Input_4(s_LOGISIM_NET_619),
                .Input_5(s_LOGISIM_NET_8),
                .Input_6(s_LOGISIM_NET_461),
                .Input_7(s_LOGISIM_NET_381),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_301),
                .Result(s_LOGISIM_NET_771));

   NOT_GATE      GATE_530 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_688));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_531 (.Input_1(s_LOGISIM_NET_131),
                .Input_2(s_LOGISIM_NET_142),
                .Input_3(s_LOGISIM_NET_402),
                .Input_4(s_LOGISIM_NET_54),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_195),
                .Input_7(s_LOGISIM_NET_354),
                .Input_8(s_LOGISIM_NET_609),
                .Result(s_LOGISIM_NET_326));

   NOT_GATE      GATE_532 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_685));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_533 (.Input_1(s_LOGISIM_NET_705),
                .Input_2(s_LOGISIM_NET_642),
                .Input_3(s_LOGISIM_NET_580),
                .Input_4(s_LOGISIM_NET_54),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_244),
                .Input_7(s_LOGISIM_NET_445),
                .Input_8(s_LOGISIM_NET_17),
                .Result(s_LOGISIM_NET_344));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_534 (.Input_1(s_LOGISIM_NET_20),
                .Input_10(s_LOGISIM_NET_159),
                .Input_2(s_LOGISIM_NET_508),
                .Input_3(s_LOGISIM_NET_7),
                .Input_4(s_LOGISIM_NET_110),
                .Input_5(s_LOGISIM_NET_8),
                .Input_6(s_LOGISIM_NET_790),
                .Input_7(s_LOGISIM_NET_430),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_80),
                .Result(s_LOGISIM_NET_493));

   NOT_GATE      GATE_535 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_34));

   NOT_GATE      GATE_536 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_617));

   NOT_GATE      GATE_537 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_108));

   NOT_GATE      GATE_538 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_135));

   NOT_GATE      GATE_539 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_479));

   NOT_GATE      GATE_540 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_627));

   NOT_GATE      GATE_541 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_708));

   NOT_GATE      GATE_542 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_206));

   NOT_GATE      GATE_543 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_294));

   NOT_GATE      GATE_544 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_419));

   NOT_GATE      GATE_545 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_274));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_546 (.Input_1(s_LOGISIM_NET_7),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_8),
                .Input_4(s_LOGISIM_NET_54),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_3),
                .Input_7(s_LOGISIM_NET_715),
                .Input_8(s_LOGISIM_NET_230),
                .Result(s_LOGISIM_NET_723));

   NOT_GATE      GATE_547 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_680));

   NOT_GATE      GATE_548 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_89));

   NOT_GATE      GATE_549 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_44));

   NOT_GATE      GATE_550 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_689));

   OR_GATE #(.BubblesMask(0))
      GATE_551 (.Input_1(s_LOGISIM_NET_484),
                .Input_2(s_LOGISIM_NET_503),
                .Result(s_LOGISIM_NET_796));

   NOT_GATE      GATE_552 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_163));

   NOT_GATE      GATE_553 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_615));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_554 (.Input_1(s_LOGISIM_NET_540),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_199),
                .Input_4(s_LOGISIM_NET_781),
                .Input_5(s_LOGISIM_NET_146),
                .Input_6(s_LOGISIM_NET_509),
                .Input_7(s_LOGISIM_NET_153),
                .Input_8(s_LOGISIM_NET_404),
                .Result(s_LOGISIM_NET_551));

   NOT_GATE      GATE_555 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_595));

   NOT_GATE      GATE_556 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_738));

   NOT_GATE      GATE_557 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_71));

   NOT_GATE      GATE_558 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_287));

   NOT_GATE      GATE_559 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_66));

   NOT_GATE      GATE_560 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_554));

   NOT_GATE      GATE_561 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_146));

   NOT_GATE      GATE_562 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_692));

   NOT_GATE      GATE_563 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_290));

   NOT_GATE      GATE_564 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_107));

   OR_GATE_29_INPUTS #(.BubblesMask(0))
      GATE_565 (.Input_1(s_LOGISIM_NET_584),
                .Input_10(s_LOGISIM_NET_379),
                .Input_11(s_LOGISIM_NET_148),
                .Input_12(s_LOGISIM_NET_389),
                .Input_13(s_LOGISIM_NET_247),
                .Input_14(s_LOGISIM_NET_493),
                .Input_15(s_LOGISIM_NET_551),
                .Input_16(s_LOGISIM_NET_378),
                .Input_17(s_LOGISIM_NET_636),
                .Input_18(s_LOGISIM_NET_326),
                .Input_19(s_LOGISIM_NET_60),
                .Input_2(s_LOGISIM_NET_338),
                .Input_20(s_LOGISIM_NET_264),
                .Input_21(s_LOGISIM_NET_697),
                .Input_22(s_LOGISIM_NET_36),
                .Input_23(s_LOGISIM_NET_255),
                .Input_24(s_LOGISIM_NET_507),
                .Input_25(s_LOGISIM_NET_481),
                .Input_26(s_LOGISIM_NET_305),
                .Input_27(s_LOGISIM_NET_176),
                .Input_28(s_LOGISIM_NET_474),
                .Input_29(s_LOGISIM_NET_563),
                .Input_3(s_LOGISIM_NET_289),
                .Input_4(s_LOGISIM_NET_0),
                .Input_5(s_LOGISIM_NET_85),
                .Input_6(s_LOGISIM_NET_756),
                .Input_7(s_LOGISIM_NET_512),
                .Input_8(s_LOGISIM_NET_316),
                .Input_9(s_LOGISIM_NET_355),
                .Result(s_LOGISIM_NET_15));

   NOT_GATE      GATE_566 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_132));

   NOT_GATE      GATE_567 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_50));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_568 (.Input_1(s_LOGISIM_NET_20),
                .Input_10(s_LOGISIM_NET_712),
                .Input_2(s_LOGISIM_NET_96),
                .Input_3(s_LOGISIM_NET_7),
                .Input_4(s_LOGISIM_NET_271),
                .Input_5(s_LOGISIM_NET_8),
                .Input_6(s_LOGISIM_NET_632),
                .Input_7(s_LOGISIM_NET_70),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_531),
                .Result(s_LOGISIM_NET_646));

   NOT_GATE      GATE_569 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_510));

   NOT_GATE      GATE_570 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_74));

   NOT_GATE      GATE_571 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_154));

   NOT_GATE      GATE_572 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_182));

   NOT_GATE      GATE_573 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_256));

   NOT_GATE      GATE_574 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_288));

   NOT_GATE      GATE_575 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_799));

   NOT_GATE      GATE_576 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_713));

   NOT_GATE      GATE_577 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_562));

   NOT_GATE      GATE_578 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_24));

   NOT_GATE      GATE_579 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_724));

   NOT_GATE      GATE_580 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_522));

   NOT_GATE      GATE_581 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_777));

   NOT_GATE      GATE_582 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_80));

   NOT_GATE      GATE_583 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_150));

   NOT_GATE      GATE_584 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_387));

   NOT_GATE      GATE_585 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_241));

   NOT_GATE      GATE_586 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_657));

   NOT_GATE      GATE_587 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_224));

   NOT_GATE      GATE_588 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_354));

   NOT_GATE      GATE_589 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_705));

   NOT_GATE      GATE_590 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_359));

   NOT_GATE      GATE_591 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_277));

   NOT_GATE      GATE_592 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_576));

   NOT_GATE      GATE_593 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_84));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_594 (.Input_1(s_LOGISIM_NET_637),
                .Input_2(s_LOGISIM_NET_576),
                .Input_3(s_LOGISIM_NET_54),
                .Input_4(s_LOGISIM_NET_287),
                .Input_5(s_LOGISIM_NET_3),
                .Input_6(s_LOGISIM_NET_349),
                .Input_7(s_LOGISIM_NET_524),
                .Result(s_LOGISIM_NET_563));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_595 (.Input_1(s_LOGISIM_NET_394),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_335),
                .Input_4(s_LOGISIM_NET_752),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_341),
                .Input_7(s_LOGISIM_NET_603),
                .Input_8(s_LOGISIM_NET_2),
                .Result(s_LOGISIM_NET_378));

   NOT_GATE      GATE_596 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_631));

   NOT_GATE      GATE_597 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_292));

   NOT_GATE      GATE_598 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_201));

   NOT_GATE      GATE_599 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_93));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_600 (.Input_1(s_LOGISIM_NET_106),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_12),
                .Input_4(s_LOGISIM_NET_672),
                .Input_5(s_LOGISIM_NET_622),
                .Input_6(s_LOGISIM_NET_29),
                .Input_7(s_LOGISIM_NET_451),
                .Input_8(s_LOGISIM_NET_667),
                .Result(s_LOGISIM_NET_484));

   NOT_GATE      GATE_601 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_11));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_602 (.Input_1(s_LOGISIM_NET_682),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_466),
                .Input_4(s_LOGISIM_NET_61),
                .Input_5(s_LOGISIM_NET_439),
                .Input_6(s_LOGISIM_NET_243),
                .Input_7(s_LOGISIM_NET_447),
                .Input_8(s_LOGISIM_NET_45),
                .Result(s_LOGISIM_NET_134));

   NOT_GATE      GATE_603 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_577));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_604 (.Input_1(s_LOGISIM_NET_242),
                .Input_2(s_LOGISIM_NET_450),
                .Input_3(s_LOGISIM_NET_54),
                .Input_4(s_LOGISIM_NET_675),
                .Input_5(s_LOGISIM_NET_3),
                .Input_6(s_LOGISIM_NET_50),
                .Input_7(s_LOGISIM_NET_459),
                .Result(s_LOGISIM_NET_467));

   NOT_GATE      GATE_605 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_579));

   NOT_GATE      GATE_606 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_156));

   NOT_GATE      GATE_607 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_227));

   NOT_GATE      GATE_608 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_518));

   NOT_GATE      GATE_609 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_785));

   NOT_GATE      GATE_610 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_696));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_611 (.Input_1(s_LOGISIM_NET_31),
                .Input_10(s_LOGISIM_NET_528),
                .Input_2(s_LOGISIM_NET_741),
                .Input_3(s_LOGISIM_NET_7),
                .Input_4(s_LOGISIM_NET_575),
                .Input_5(s_LOGISIM_NET_8),
                .Input_6(s_LOGISIM_NET_398),
                .Input_7(s_LOGISIM_NET_291),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_200),
                .Result(s_LOGISIM_NET_332));

   NOT_GATE      GATE_612 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_366));

   NOT_GATE      GATE_613 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_504));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_614 (.Input_1(s_LOGISIM_NET_172),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_312),
                .Input_4(s_LOGISIM_NET_601),
                .Input_5(s_LOGISIM_NET_541),
                .Input_6(s_LOGISIM_NET_139),
                .Input_7(s_LOGISIM_NET_327),
                .Input_8(s_LOGISIM_NET_596),
                .Result(s_LOGISIM_NET_598));

   NOT_GATE      GATE_615 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_151));

   OR_GATE_3_INPUTS #(.BubblesMask(0))
      GATE_616 (.Input_1(s_LOGISIM_NET_165),
                .Input_2(s_LOGISIM_NET_797),
                .Input_3(s_LOGISIM_NET_436),
                .Result(s_LOGISIM_NET_778));

   NOT_GATE      GATE_617 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_314));

   NOT_GATE      GATE_618 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_681));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_619 (.Input_1(s_LOGISIM_NET_240),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_152),
                .Input_4(s_LOGISIM_NET_704),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_166),
                .Input_7(s_LOGISIM_NET_518),
                .Input_8(s_LOGISIM_NET_17),
                .Result(s_LOGISIM_NET_683));

   NOT_GATE      GATE_620 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_315));

   NOT_GATE      GATE_621 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_444));

   NOT_GATE      GATE_622 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_499));

   NOT_GATE      GATE_623 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_677));

   NOT_GATE      GATE_624 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_573));

   NOT_GATE      GATE_625 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_525));

   NOT_GATE      GATE_626 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_130));

   NOT_GATE      GATE_627 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_244));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_628 (.Input_1(s_LOGISIM_NET_497),
                .Input_10(s_LOGISIM_NET_788),
                .Input_2(s_LOGISIM_NET_431),
                .Input_3(s_LOGISIM_NET_7),
                .Input_4(s_LOGISIM_NET_9),
                .Input_5(s_LOGISIM_NET_8),
                .Input_6(s_LOGISIM_NET_760),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_717),
                .Result(s_LOGISIM_NET_289));

   NOT_GATE      GATE_629 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_618));

   NOT_GATE      GATE_630 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_249));

   NOT_GATE      GATE_631 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_721));

   NOT_GATE      GATE_632 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_114));

   NOT_GATE      GATE_633 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_625));

   NOT_GATE      GATE_634 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_655));

   NOT_GATE      GATE_635 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_578));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_636 (.Input_1(s_LOGISIM_NET_44),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_224),
                .Input_4(s_LOGISIM_NET_558),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_13),
                .Input_7(s_LOGISIM_NET_238),
                .Input_8(s_LOGISIM_NET_17),
                .Result(s_LOGISIM_NET_122));

   NOT_GATE      GATE_637 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_167));

   NOT_GATE      GATE_638 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_454));

   NOT_GATE      GATE_639 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_649));

   NOT_GATE      GATE_640 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_222));

   NOT_GATE      GATE_641 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_331));

   NOT_GATE      GATE_642 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_377));

   AND_GATE_5_INPUTS #(.BubblesMask(0))
      GATE_643 (.Input_1(s_LOGISIM_NET_182),
                .Input_2(s_LOGISIM_NET_21),
                .Input_3(s_LOGISIM_NET_3),
                .Input_4(s_LOGISIM_NET_56),
                .Input_5(s_LOGISIM_NET_17),
                .Result(s_LOGISIM_NET_190));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_644 (.Input_1(s_LOGISIM_NET_7),
                .Input_2(s_LOGISIM_NET_695),
                .Input_3(s_LOGISIM_NET_8),
                .Input_4(s_LOGISIM_NET_294),
                .Input_5(s_LOGISIM_NET_158),
                .Input_6(s_LOGISIM_NET_407),
                .Input_7(s_LOGISIM_NET_568),
                .Input_8(s_LOGISIM_NET_288),
                .Result(s_LOGISIM_NET_791));

   NOT_GATE      GATE_645 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_157));

   NOT_GATE      GATE_646 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_217));

   NOT_GATE      GATE_647 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_453));

   NOT_GATE      GATE_648 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_714));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_649 (.Input_1(s_LOGISIM_NET_20),
                .Input_10(s_LOGISIM_NET_773),
                .Input_2(s_LOGISIM_NET_261),
                .Input_3(s_LOGISIM_NET_377),
                .Input_4(s_LOGISIM_NET_147),
                .Input_5(s_LOGISIM_NET_708),
                .Input_6(s_LOGISIM_NET_24),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_676),
                .Result(s_LOGISIM_NET_358));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_650 (.Input_1(s_LOGISIM_NET_20),
                .Input_10(s_LOGISIM_NET_371),
                .Input_2(s_LOGISIM_NET_664),
                .Input_3(s_LOGISIM_NET_7),
                .Input_4(s_LOGISIM_NET_427),
                .Input_5(s_LOGISIM_NET_8),
                .Input_6(s_LOGISIM_NET_163),
                .Input_7(s_LOGISIM_NET_613),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_123),
                .Result(s_LOGISIM_NET_38));

   NOT_GATE      GATE_651 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_166));

   NOT_GATE      GATE_652 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_744));

   NOT_GATE      GATE_653 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_168));

   NOT_GATE      GATE_654 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_559));

   NOT_GATE      GATE_655 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_72));

   NOT_GATE      GATE_656 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_605));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_657 (.Input_1(s_LOGISIM_NET_256),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_174),
                .Input_4(s_LOGISIM_NET_711),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_188),
                .Input_7(s_LOGISIM_NET_523),
                .Input_8(s_LOGISIM_NET_17),
                .Result(s_LOGISIM_NET_176));

   NOT_GATE      GATE_658 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_271));

   NOT_GATE      GATE_659 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_533));

   NOT_GATE      GATE_660 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_754));

   NOT_GATE      GATE_661 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_46));

   NOT_GATE      GATE_662 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_491));

   NOT_GATE      GATE_663 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_195));

   NOT_GATE      GATE_664 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_541));

   NOT_GATE      GATE_665 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_545));

   NOT_GATE      GATE_666 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_488));

   NOT_GATE      GATE_667 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_109));

   NOT_GATE      GATE_668 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_735));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_669 (.Input_1(s_LOGISIM_NET_292),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_221),
                .Input_4(s_LOGISIM_NET_721),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_232),
                .Input_7(s_LOGISIM_NET_546),
                .Input_8(s_LOGISIM_NET_17),
                .Result(s_LOGISIM_NET_663));

   NOT_GATE      GATE_670 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_515));

   NOT_GATE      GATE_671 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_81));

   NOT_GATE      GATE_672 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_568));

   NOT_GATE      GATE_673 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_675));

   NOT_GATE      GATE_674 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_539));

   NOT_GATE      GATE_675 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_279));

   NOT_GATE      GATE_676 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_693));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_677 (.Input_1(s_LOGISIM_NET_599),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_310),
                .Input_4(s_LOGISIM_NET_792),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_573),
                .Input_7(s_LOGISIM_NET_136),
                .Input_8(s_LOGISIM_NET_17),
                .Result(s_LOGISIM_NET_740));

   NOT_GATE      GATE_678 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_616));

   NOT_GATE      GATE_679 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_343));

   NOT_GATE      GATE_680 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_779));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_681 (.Input_1(s_LOGISIM_NET_729),
                .Input_10(s_LOGISIM_NET_449),
                .Input_2(s_LOGISIM_NET_701),
                .Input_3(s_LOGISIM_NET_641),
                .Input_4(s_LOGISIM_NET_9),
                .Input_5(s_LOGISIM_NET_8),
                .Input_6(s_LOGISIM_NET_297),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_28),
                .Result(s_LOGISIM_NET_88));

   OR_GATE #(.BubblesMask(0))
      GATE_682 (.Input_1(s_LOGISIM_NET_467),
                .Input_2(s_LOGISIM_NET_121),
                .Result(s_LOGISIM_NET_728));

   NOT_GATE      GATE_683 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_64));

   NOT_GATE      GATE_684 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_653));

   NOT_GATE      GATE_685 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_425));

   NOT_GATE      GATE_686 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_581));

   NOT_GATE      GATE_687 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_582));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_688 (.Input_1(s_LOGISIM_NET_233),
                .Input_10(s_LOGISIM_NET_6),
                .Input_2(s_LOGISIM_NET_128),
                .Input_3(s_LOGISIM_NET_443),
                .Input_4(s_LOGISIM_NET_279),
                .Input_5(s_LOGISIM_NET_737),
                .Input_6(s_LOGISIM_NET_169),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_713),
                .Result(s_LOGISIM_NET_105));

   NOT_GATE      GATE_689 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_252));

   NOT_GATE      GATE_690 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_14));

   NOT_GATE      GATE_691 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_236));

   NOT_GATE      GATE_692 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_262));

   NOT_GATE      GATE_693 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_684));

   NOT_GATE      GATE_694 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_502));

   NOT_GATE      GATE_695 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_706));

   NOT_GATE      GATE_696 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_173));

   NOT_GATE      GATE_697 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_556));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_698 (.Input_1(s_LOGISIM_NET_246),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_156),
                .Input_4(s_LOGISIM_NET_707),
                .Input_5(s_LOGISIM_NET_22),
                .Input_6(s_LOGISIM_NET_177),
                .Input_7(s_LOGISIM_NET_522),
                .Input_8(s_LOGISIM_NET_17),
                .Result(s_LOGISIM_NET_762));

   NOT_GATE      GATE_699 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_731));

   NOT_GATE      GATE_700 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_594));

   NOT_GATE      GATE_701 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_320));

   NOT_GATE      GATE_702 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_764));

   NOT_GATE      GATE_703 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_586));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_704 (.Input_1(s_LOGISIM_NET_7),
                .Input_2(s_LOGISIM_NET_359),
                .Input_3(s_LOGISIM_NET_8),
                .Input_4(s_LOGISIM_NET_696),
                .Input_5(s_LOGISIM_NET_653),
                .Input_6(s_LOGISIM_NET_135),
                .Input_7(s_LOGISIM_NET_505),
                .Input_8(s_LOGISIM_NET_693),
                .Result(s_LOGISIM_NET_36));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_705 (.Input_1(s_LOGISIM_NET_83),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_257),
                .Input_4(s_LOGISIM_NET_572),
                .Input_5(s_LOGISIM_NET_504),
                .Input_6(s_LOGISIM_NET_52),
                .Input_7(s_LOGISIM_NET_276),
                .Input_8(s_LOGISIM_NET_17),
                .Result(s_LOGISIM_NET_503));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_706 (.Input_1(s_LOGISIM_NET_7),
                .Input_2(s_LOGISIM_NET_700),
                .Input_3(s_LOGISIM_NET_8),
                .Input_4(s_LOGISIM_NET_54),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_274),
                .Input_7(s_LOGISIM_NET_463),
                .Input_8(s_LOGISIM_NET_249),
                .Result(s_LOGISIM_NET_309));

   NOT_GATE      GATE_707 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_169));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_708 (.Input_1(s_LOGISIM_NET_206),
                .Input_10(s_LOGISIM_NET_749),
                .Input_2(s_LOGISIM_NET_87),
                .Input_3(s_LOGISIM_NET_7),
                .Input_4(s_LOGISIM_NET_9),
                .Input_5(s_LOGISIM_NET_635),
                .Input_6(s_LOGISIM_NET_557),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_602),
                .Result(s_LOGISIM_NET_0));

   NOT_GATE      GATE_709 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_349));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_710 (.Input_1(s_LOGISIM_NET_7),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_308),
                .Input_4(s_LOGISIM_NET_745),
                .Input_5(s_LOGISIM_NET_217),
                .Input_6(s_LOGISIM_NET_3),
                .Input_7(s_LOGISIM_NET_588),
                .Input_8(s_LOGISIM_NET_743),
                .Result(s_LOGISIM_NET_355));

   NOT_GATE      GATE_711 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_348));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_712 (.Input_1(s_LOGISIM_NET_699),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_502),
                .Input_4(s_LOGISIM_NET_129),
                .Input_5(s_LOGISIM_NET_478),
                .Input_6(s_LOGISIM_NET_293),
                .Input_7(s_LOGISIM_NET_480),
                .Input_8(s_LOGISIM_NET_17),
                .Result(s_LOGISIM_NET_42));

   NOT_GATE      GATE_713 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_199));

   NOT_GATE      GATE_714 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_790));

   NOT_GATE      GATE_715 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_709));

   NOT_GATE      GATE_716 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_786));

   NOT_GATE      GATE_717 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_800));

   NOT_GATE      GATE_718 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_398));

   NOT_GATE      GATE_719 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_393));

   NOT_GATE      GATE_720 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_606));

   NOT_GATE      GATE_721 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_381));

   NOT_GATE      GATE_722 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_162));

   NOT_GATE      GATE_723 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_164));

   NOT_GATE      GATE_724 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_302));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_725 (.Input_1(s_LOGISIM_NET_250),
                .Input_2(s_LOGISIM_NET_311),
                .Input_3(s_LOGISIM_NET_53),
                .Input_4(s_LOGISIM_NET_679),
                .Input_5(s_LOGISIM_NET_629),
                .Input_6(s_LOGISIM_NET_3),
                .Input_7(s_LOGISIM_NET_465),
                .Input_8(s_LOGISIM_NET_673),
                .Result(s_LOGISIM_NET_726));

   NOT_GATE      GATE_726 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_94));

   NOT_GATE      GATE_727 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_179));

   NOT_GATE      GATE_728 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_126));

   NOT_GATE      GATE_729 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_365));

   NOT_GATE      GATE_730 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_652));

   NOT_GATE      GATE_731 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_321));

   NOT_GATE      GATE_732 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_276));

   NOT_GATE      GATE_733 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_386));

   NOT_GATE      GATE_734 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_715));

   NOT_GATE      GATE_735 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_188));

   NOT_GATE      GATE_736 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_212));

   NOT_GATE      GATE_737 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_789));

   NOT_GATE      GATE_738 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_323));

   NOT_GATE      GATE_739 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_475));

   NOT_GATE      GATE_740 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_284));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_741 (.Input_1(s_LOGISIM_NET_628),
                .Input_2(s_LOGISIM_NET_555),
                .Input_3(s_LOGISIM_NET_54),
                .Input_4(s_LOGISIM_NET_251),
                .Input_5(s_LOGISIM_NET_3),
                .Input_6(s_LOGISIM_NET_313),
                .Input_7(s_LOGISIM_NET_501),
                .Result(s_LOGISIM_NET_18));

   NOT_GATE      GATE_742 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_420));

   NOT_GATE      GATE_743 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_798));

   NOT_GATE      GATE_744 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_619));

   NOT_GATE      GATE_745 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_793));

   NOT_GATE      GATE_746 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_639));

   NOT_GATE      GATE_747 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_775));

   NOT_GATE      GATE_748 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_628));

   NOT_GATE      GATE_749 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_189));

   NOT_GATE      GATE_750 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_317));

   NOT_GATE      GATE_751 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_295));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_752 (.Input_1(s_LOGISIM_NET_462),
                .Input_10(s_LOGISIM_NET_47),
                .Input_2(s_LOGISIM_NET_409),
                .Input_3(s_LOGISIM_NET_283),
                .Input_4(s_LOGISIM_NET_86),
                .Input_5(s_LOGISIM_NET_779),
                .Input_6(s_LOGISIM_NET_54),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_3),
                .Input_9(s_LOGISIM_NET_767),
                .Result(s_LOGISIM_NET_514));

   NOT_GATE      GATE_753 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_700));

   NOT_GATE      GATE_754 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_674));

   NOT_GATE      GATE_755 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_124));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_756 (.Input_1(s_LOGISIM_NET_543),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_193),
                .Input_4(s_LOGISIM_NET_783),
                .Input_5(s_LOGISIM_NET_151),
                .Input_6(s_LOGISIM_NET_3),
                .Input_7(s_LOGISIM_NET_694),
                .Input_8(s_LOGISIM_NET_300),
                .Result(s_LOGISIM_NET_725));

   NOT_GATE      GATE_757 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_801));

   NOT_GATE      GATE_758 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_293));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_759 (.Input_1(s_LOGISIM_NET_630),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_376),
                .Input_4(s_LOGISIM_NET_801),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_608),
                .Input_7(s_LOGISIM_NET_239),
                .Input_8(s_LOGISIM_NET_17),
                .Result(s_LOGISIM_NET_794));

   NOT_GATE      GATE_760 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_258));

   NOT_GATE      GATE_761 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_102));

   NOT_GATE      GATE_762 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_470));

   NOT_GATE      GATE_763 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_621));

   NOT_GATE      GATE_764 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_73));

   NOT_GATE      GATE_765 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_783));

   NOT_GATE      GATE_766 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_137));

   OR_GATE_4_INPUTS #(.BubblesMask(0))
      GATE_767 (.Input_1(s_LOGISIM_NET_145),
                .Input_2(s_LOGISIM_NET_372),
                .Input_3(s_LOGISIM_NET_18),
                .Input_4(s_LOGISIM_NET_339),
                .Result(s_LOGISIM_NET_736));

   NOT_GATE      GATE_768 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_383));

   NOT_GATE      GATE_769 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_191));

   NOT_GATE      GATE_770 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_613));

   NOT_GATE      GATE_771 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_406));

   NOT_GATE      GATE_772 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_342));

   NOT_GATE      GATE_773 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_62));

   NOT_GATE      GATE_774 (.Input_1(s_LOGISIM_NET_8),
                           .Result(s_LOGISIM_NET_537));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_775 (.Input_1(s_LOGISIM_NET_684),
                .Input_2(s_LOGISIM_NET_620),
                .Input_3(s_LOGISIM_NET_54),
                .Input_4(s_LOGISIM_NET_375),
                .Input_5(s_LOGISIM_NET_3),
                .Input_6(s_LOGISIM_NET_423),
                .Input_7(s_LOGISIM_NET_14),
                .Result(s_LOGISIM_NET_121));

   NOT_GATE      GATE_776 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_334));

   NOT_GATE      GATE_777 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_83));

   NOT_GATE      GATE_778 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_449));

   NOT_GATE      GATE_779 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_459));

   NOT_GATE      GATE_780 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_43));

   NOT_GATE      GATE_781 (.Input_1(s_LOGISIM_NET_20),
                           .Result(s_LOGISIM_NET_265));

   NOT_GATE      GATE_782 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_534));

   NOT_GATE      GATE_783 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_370));

   NOT_GATE      GATE_784 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_717));

   NOT_GATE      GATE_785 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_118));

   NOT_GATE      GATE_786 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_418));

   NOT_GATE      GATE_787 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_429));

   NOT_GATE      GATE_788 (.Input_1(s_LOGISIM_NET_54),
                           .Result(s_LOGISIM_NET_760));

   NOT_GATE      GATE_789 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_440));

   NOT_GATE      GATE_790 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_161));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_791 (.Input_1(s_LOGISIM_NET_678),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_456),
                .Input_4(s_LOGISIM_NET_39),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_58),
                .Input_7(s_LOGISIM_NET_347),
                .Input_8(s_LOGISIM_NET_19),
                .Result(s_LOGISIM_NET_37));

   NOT_GATE      GATE_792 (.Input_1(s_LOGISIM_NET_21),
                           .Result(s_LOGISIM_NET_333));

   NOT_GATE      GATE_793 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_139));

   NOT_GATE      GATE_794 (.Input_1(s_LOGISIM_NET_17),
                           .Result(s_LOGISIM_NET_437));

   NOT_GATE      GATE_795 (.Input_1(s_LOGISIM_NET_3),
                           .Result(s_LOGISIM_NET_207));



endmodule
